// test

module \AND2  ( 
    \V1 , \V2 ,
    \W1 );
  input  \V1 , \V2 ;
  output \W1 ;
  
  assign \W1 = \V1 & \V2  ;
endmodule


