// Benchmark "Sorter100" written by ABC on Tue Apr  9 09:15:00 2024

module Sorter100 ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27,
    x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41,
    x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55,
    x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69,
    x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83,
    x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97,
    x98, x99,
    y00, y01, y02, y03, y04, y05, y06, y07, y08, y09, y10, y11, y12, y13,
    y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27,
    y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41,
    y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55,
    y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69,
    y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83,
    y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97,
    y98, y99  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26,
    x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40,
    x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54,
    x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68,
    x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82,
    x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96,
    x97, x98, x99;
  output y00, y01, y02, y03, y04, y05, y06, y07, y08, y09, y10, y11, y12, y13,
    y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27,
    y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41,
    y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55,
    y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69,
    y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83,
    y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97,
    y98, y99;
  wire \new_Sorter100|0000_ , \new_Sorter100|0001_ , \new_Sorter100|0002_ ,
    \new_Sorter100|0003_ , \new_Sorter100|0004_ , \new_Sorter100|0005_ ,
    \new_Sorter100|0006_ , \new_Sorter100|0007_ , \new_Sorter100|0008_ ,
    \new_Sorter100|0009_ , \new_Sorter100|0010_ , \new_Sorter100|0011_ ,
    \new_Sorter100|0012_ , \new_Sorter100|0013_ , \new_Sorter100|0014_ ,
    \new_Sorter100|0015_ , \new_Sorter100|0016_ , \new_Sorter100|0017_ ,
    \new_Sorter100|0018_ , \new_Sorter100|0019_ , \new_Sorter100|0020_ ,
    \new_Sorter100|0021_ , \new_Sorter100|0022_ , \new_Sorter100|0023_ ,
    \new_Sorter100|0024_ , \new_Sorter100|0025_ , \new_Sorter100|0026_ ,
    \new_Sorter100|0027_ , \new_Sorter100|0028_ , \new_Sorter100|0029_ ,
    \new_Sorter100|0030_ , \new_Sorter100|0031_ , \new_Sorter100|0032_ ,
    \new_Sorter100|0033_ , \new_Sorter100|0034_ , \new_Sorter100|0035_ ,
    \new_Sorter100|0036_ , \new_Sorter100|0037_ , \new_Sorter100|0038_ ,
    \new_Sorter100|0039_ , \new_Sorter100|0040_ , \new_Sorter100|0041_ ,
    \new_Sorter100|0042_ , \new_Sorter100|0043_ , \new_Sorter100|0044_ ,
    \new_Sorter100|0045_ , \new_Sorter100|0046_ , \new_Sorter100|0047_ ,
    \new_Sorter100|0048_ , \new_Sorter100|0049_ , \new_Sorter100|0050_ ,
    \new_Sorter100|0051_ , \new_Sorter100|0052_ , \new_Sorter100|0053_ ,
    \new_Sorter100|0054_ , \new_Sorter100|0055_ , \new_Sorter100|0056_ ,
    \new_Sorter100|0057_ , \new_Sorter100|0058_ , \new_Sorter100|0059_ ,
    \new_Sorter100|0060_ , \new_Sorter100|0061_ , \new_Sorter100|0062_ ,
    \new_Sorter100|0063_ , \new_Sorter100|0064_ , \new_Sorter100|0065_ ,
    \new_Sorter100|0066_ , \new_Sorter100|0067_ , \new_Sorter100|0068_ ,
    \new_Sorter100|0069_ , \new_Sorter100|0070_ , \new_Sorter100|0071_ ,
    \new_Sorter100|0072_ , \new_Sorter100|0073_ , \new_Sorter100|0074_ ,
    \new_Sorter100|0075_ , \new_Sorter100|0076_ , \new_Sorter100|0077_ ,
    \new_Sorter100|0078_ , \new_Sorter100|0079_ , \new_Sorter100|0080_ ,
    \new_Sorter100|0081_ , \new_Sorter100|0082_ , \new_Sorter100|0083_ ,
    \new_Sorter100|0084_ , \new_Sorter100|0085_ , \new_Sorter100|0086_ ,
    \new_Sorter100|0087_ , \new_Sorter100|0088_ , \new_Sorter100|0089_ ,
    \new_Sorter100|0090_ , \new_Sorter100|0091_ , \new_Sorter100|0092_ ,
    \new_Sorter100|0093_ , \new_Sorter100|0094_ , \new_Sorter100|0095_ ,
    \new_Sorter100|0096_ , \new_Sorter100|0097_ , \new_Sorter100|0098_ ,
    \new_Sorter100|0099_ , \new_Sorter100|0100_ , \new_Sorter100|0199_ ,
    \new_Sorter100|0101_ , \new_Sorter100|0102_ , \new_Sorter100|0103_ ,
    \new_Sorter100|0104_ , \new_Sorter100|0105_ , \new_Sorter100|0106_ ,
    \new_Sorter100|0107_ , \new_Sorter100|0108_ , \new_Sorter100|0109_ ,
    \new_Sorter100|0110_ , \new_Sorter100|0111_ , \new_Sorter100|0112_ ,
    \new_Sorter100|0113_ , \new_Sorter100|0114_ , \new_Sorter100|0115_ ,
    \new_Sorter100|0116_ , \new_Sorter100|0117_ , \new_Sorter100|0118_ ,
    \new_Sorter100|0119_ , \new_Sorter100|0120_ , \new_Sorter100|0121_ ,
    \new_Sorter100|0122_ , \new_Sorter100|0123_ , \new_Sorter100|0124_ ,
    \new_Sorter100|0125_ , \new_Sorter100|0126_ , \new_Sorter100|0127_ ,
    \new_Sorter100|0128_ , \new_Sorter100|0129_ , \new_Sorter100|0130_ ,
    \new_Sorter100|0131_ , \new_Sorter100|0132_ , \new_Sorter100|0133_ ,
    \new_Sorter100|0134_ , \new_Sorter100|0135_ , \new_Sorter100|0136_ ,
    \new_Sorter100|0137_ , \new_Sorter100|0138_ , \new_Sorter100|0139_ ,
    \new_Sorter100|0140_ , \new_Sorter100|0141_ , \new_Sorter100|0142_ ,
    \new_Sorter100|0143_ , \new_Sorter100|0144_ , \new_Sorter100|0145_ ,
    \new_Sorter100|0146_ , \new_Sorter100|0147_ , \new_Sorter100|0148_ ,
    \new_Sorter100|0149_ , \new_Sorter100|0150_ , \new_Sorter100|0151_ ,
    \new_Sorter100|0152_ , \new_Sorter100|0153_ , \new_Sorter100|0154_ ,
    \new_Sorter100|0155_ , \new_Sorter100|0156_ , \new_Sorter100|0157_ ,
    \new_Sorter100|0158_ , \new_Sorter100|0159_ , \new_Sorter100|0160_ ,
    \new_Sorter100|0161_ , \new_Sorter100|0162_ , \new_Sorter100|0163_ ,
    \new_Sorter100|0164_ , \new_Sorter100|0165_ , \new_Sorter100|0166_ ,
    \new_Sorter100|0167_ , \new_Sorter100|0168_ , \new_Sorter100|0169_ ,
    \new_Sorter100|0170_ , \new_Sorter100|0171_ , \new_Sorter100|0172_ ,
    \new_Sorter100|0173_ , \new_Sorter100|0174_ , \new_Sorter100|0175_ ,
    \new_Sorter100|0176_ , \new_Sorter100|0177_ , \new_Sorter100|0178_ ,
    \new_Sorter100|0179_ , \new_Sorter100|0180_ , \new_Sorter100|0181_ ,
    \new_Sorter100|0182_ , \new_Sorter100|0183_ , \new_Sorter100|0184_ ,
    \new_Sorter100|0185_ , \new_Sorter100|0186_ , \new_Sorter100|0187_ ,
    \new_Sorter100|0188_ , \new_Sorter100|0189_ , \new_Sorter100|0190_ ,
    \new_Sorter100|0191_ , \new_Sorter100|0192_ , \new_Sorter100|0193_ ,
    \new_Sorter100|0194_ , \new_Sorter100|0195_ , \new_Sorter100|0196_ ,
    \new_Sorter100|0197_ , \new_Sorter100|0198_ , \new_Sorter100|0200_ ,
    \new_Sorter100|0201_ , \new_Sorter100|0202_ , \new_Sorter100|0203_ ,
    \new_Sorter100|0204_ , \new_Sorter100|0205_ , \new_Sorter100|0206_ ,
    \new_Sorter100|0207_ , \new_Sorter100|0208_ , \new_Sorter100|0209_ ,
    \new_Sorter100|0210_ , \new_Sorter100|0211_ , \new_Sorter100|0212_ ,
    \new_Sorter100|0213_ , \new_Sorter100|0214_ , \new_Sorter100|0215_ ,
    \new_Sorter100|0216_ , \new_Sorter100|0217_ , \new_Sorter100|0218_ ,
    \new_Sorter100|0219_ , \new_Sorter100|0220_ , \new_Sorter100|0221_ ,
    \new_Sorter100|0222_ , \new_Sorter100|0223_ , \new_Sorter100|0224_ ,
    \new_Sorter100|0225_ , \new_Sorter100|0226_ , \new_Sorter100|0227_ ,
    \new_Sorter100|0228_ , \new_Sorter100|0229_ , \new_Sorter100|0230_ ,
    \new_Sorter100|0231_ , \new_Sorter100|0232_ , \new_Sorter100|0233_ ,
    \new_Sorter100|0234_ , \new_Sorter100|0235_ , \new_Sorter100|0236_ ,
    \new_Sorter100|0237_ , \new_Sorter100|0238_ , \new_Sorter100|0239_ ,
    \new_Sorter100|0240_ , \new_Sorter100|0241_ , \new_Sorter100|0242_ ,
    \new_Sorter100|0243_ , \new_Sorter100|0244_ , \new_Sorter100|0245_ ,
    \new_Sorter100|0246_ , \new_Sorter100|0247_ , \new_Sorter100|0248_ ,
    \new_Sorter100|0249_ , \new_Sorter100|0250_ , \new_Sorter100|0251_ ,
    \new_Sorter100|0252_ , \new_Sorter100|0253_ , \new_Sorter100|0254_ ,
    \new_Sorter100|0255_ , \new_Sorter100|0256_ , \new_Sorter100|0257_ ,
    \new_Sorter100|0258_ , \new_Sorter100|0259_ , \new_Sorter100|0260_ ,
    \new_Sorter100|0261_ , \new_Sorter100|0262_ , \new_Sorter100|0263_ ,
    \new_Sorter100|0264_ , \new_Sorter100|0265_ , \new_Sorter100|0266_ ,
    \new_Sorter100|0267_ , \new_Sorter100|0268_ , \new_Sorter100|0269_ ,
    \new_Sorter100|0270_ , \new_Sorter100|0271_ , \new_Sorter100|0272_ ,
    \new_Sorter100|0273_ , \new_Sorter100|0274_ , \new_Sorter100|0275_ ,
    \new_Sorter100|0276_ , \new_Sorter100|0277_ , \new_Sorter100|0278_ ,
    \new_Sorter100|0279_ , \new_Sorter100|0280_ , \new_Sorter100|0281_ ,
    \new_Sorter100|0282_ , \new_Sorter100|0283_ , \new_Sorter100|0284_ ,
    \new_Sorter100|0285_ , \new_Sorter100|0286_ , \new_Sorter100|0287_ ,
    \new_Sorter100|0288_ , \new_Sorter100|0289_ , \new_Sorter100|0290_ ,
    \new_Sorter100|0291_ , \new_Sorter100|0292_ , \new_Sorter100|0293_ ,
    \new_Sorter100|0294_ , \new_Sorter100|0295_ , \new_Sorter100|0296_ ,
    \new_Sorter100|0297_ , \new_Sorter100|0298_ , \new_Sorter100|0299_ ,
    \new_Sorter100|0300_ , \new_Sorter100|0399_ , \new_Sorter100|0301_ ,
    \new_Sorter100|0302_ , \new_Sorter100|0303_ , \new_Sorter100|0304_ ,
    \new_Sorter100|0305_ , \new_Sorter100|0306_ , \new_Sorter100|0307_ ,
    \new_Sorter100|0308_ , \new_Sorter100|0309_ , \new_Sorter100|0310_ ,
    \new_Sorter100|0311_ , \new_Sorter100|0312_ , \new_Sorter100|0313_ ,
    \new_Sorter100|0314_ , \new_Sorter100|0315_ , \new_Sorter100|0316_ ,
    \new_Sorter100|0317_ , \new_Sorter100|0318_ , \new_Sorter100|0319_ ,
    \new_Sorter100|0320_ , \new_Sorter100|0321_ , \new_Sorter100|0322_ ,
    \new_Sorter100|0323_ , \new_Sorter100|0324_ , \new_Sorter100|0325_ ,
    \new_Sorter100|0326_ , \new_Sorter100|0327_ , \new_Sorter100|0328_ ,
    \new_Sorter100|0329_ , \new_Sorter100|0330_ , \new_Sorter100|0331_ ,
    \new_Sorter100|0332_ , \new_Sorter100|0333_ , \new_Sorter100|0334_ ,
    \new_Sorter100|0335_ , \new_Sorter100|0336_ , \new_Sorter100|0337_ ,
    \new_Sorter100|0338_ , \new_Sorter100|0339_ , \new_Sorter100|0340_ ,
    \new_Sorter100|0341_ , \new_Sorter100|0342_ , \new_Sorter100|0343_ ,
    \new_Sorter100|0344_ , \new_Sorter100|0345_ , \new_Sorter100|0346_ ,
    \new_Sorter100|0347_ , \new_Sorter100|0348_ , \new_Sorter100|0349_ ,
    \new_Sorter100|0350_ , \new_Sorter100|0351_ , \new_Sorter100|0352_ ,
    \new_Sorter100|0353_ , \new_Sorter100|0354_ , \new_Sorter100|0355_ ,
    \new_Sorter100|0356_ , \new_Sorter100|0357_ , \new_Sorter100|0358_ ,
    \new_Sorter100|0359_ , \new_Sorter100|0360_ , \new_Sorter100|0361_ ,
    \new_Sorter100|0362_ , \new_Sorter100|0363_ , \new_Sorter100|0364_ ,
    \new_Sorter100|0365_ , \new_Sorter100|0366_ , \new_Sorter100|0367_ ,
    \new_Sorter100|0368_ , \new_Sorter100|0369_ , \new_Sorter100|0370_ ,
    \new_Sorter100|0371_ , \new_Sorter100|0372_ , \new_Sorter100|0373_ ,
    \new_Sorter100|0374_ , \new_Sorter100|0375_ , \new_Sorter100|0376_ ,
    \new_Sorter100|0377_ , \new_Sorter100|0378_ , \new_Sorter100|0379_ ,
    \new_Sorter100|0380_ , \new_Sorter100|0381_ , \new_Sorter100|0382_ ,
    \new_Sorter100|0383_ , \new_Sorter100|0384_ , \new_Sorter100|0385_ ,
    \new_Sorter100|0386_ , \new_Sorter100|0387_ , \new_Sorter100|0388_ ,
    \new_Sorter100|0389_ , \new_Sorter100|0390_ , \new_Sorter100|0391_ ,
    \new_Sorter100|0392_ , \new_Sorter100|0393_ , \new_Sorter100|0394_ ,
    \new_Sorter100|0395_ , \new_Sorter100|0396_ , \new_Sorter100|0397_ ,
    \new_Sorter100|0398_ , \new_Sorter100|0400_ , \new_Sorter100|0401_ ,
    \new_Sorter100|0402_ , \new_Sorter100|0403_ , \new_Sorter100|0404_ ,
    \new_Sorter100|0405_ , \new_Sorter100|0406_ , \new_Sorter100|0407_ ,
    \new_Sorter100|0408_ , \new_Sorter100|0409_ , \new_Sorter100|0410_ ,
    \new_Sorter100|0411_ , \new_Sorter100|0412_ , \new_Sorter100|0413_ ,
    \new_Sorter100|0414_ , \new_Sorter100|0415_ , \new_Sorter100|0416_ ,
    \new_Sorter100|0417_ , \new_Sorter100|0418_ , \new_Sorter100|0419_ ,
    \new_Sorter100|0420_ , \new_Sorter100|0421_ , \new_Sorter100|0422_ ,
    \new_Sorter100|0423_ , \new_Sorter100|0424_ , \new_Sorter100|0425_ ,
    \new_Sorter100|0426_ , \new_Sorter100|0427_ , \new_Sorter100|0428_ ,
    \new_Sorter100|0429_ , \new_Sorter100|0430_ , \new_Sorter100|0431_ ,
    \new_Sorter100|0432_ , \new_Sorter100|0433_ , \new_Sorter100|0434_ ,
    \new_Sorter100|0435_ , \new_Sorter100|0436_ , \new_Sorter100|0437_ ,
    \new_Sorter100|0438_ , \new_Sorter100|0439_ , \new_Sorter100|0440_ ,
    \new_Sorter100|0441_ , \new_Sorter100|0442_ , \new_Sorter100|0443_ ,
    \new_Sorter100|0444_ , \new_Sorter100|0445_ , \new_Sorter100|0446_ ,
    \new_Sorter100|0447_ , \new_Sorter100|0448_ , \new_Sorter100|0449_ ,
    \new_Sorter100|0450_ , \new_Sorter100|0451_ , \new_Sorter100|0452_ ,
    \new_Sorter100|0453_ , \new_Sorter100|0454_ , \new_Sorter100|0455_ ,
    \new_Sorter100|0456_ , \new_Sorter100|0457_ , \new_Sorter100|0458_ ,
    \new_Sorter100|0459_ , \new_Sorter100|0460_ , \new_Sorter100|0461_ ,
    \new_Sorter100|0462_ , \new_Sorter100|0463_ , \new_Sorter100|0464_ ,
    \new_Sorter100|0465_ , \new_Sorter100|0466_ , \new_Sorter100|0467_ ,
    \new_Sorter100|0468_ , \new_Sorter100|0469_ , \new_Sorter100|0470_ ,
    \new_Sorter100|0471_ , \new_Sorter100|0472_ , \new_Sorter100|0473_ ,
    \new_Sorter100|0474_ , \new_Sorter100|0475_ , \new_Sorter100|0476_ ,
    \new_Sorter100|0477_ , \new_Sorter100|0478_ , \new_Sorter100|0479_ ,
    \new_Sorter100|0480_ , \new_Sorter100|0481_ , \new_Sorter100|0482_ ,
    \new_Sorter100|0483_ , \new_Sorter100|0484_ , \new_Sorter100|0485_ ,
    \new_Sorter100|0486_ , \new_Sorter100|0487_ , \new_Sorter100|0488_ ,
    \new_Sorter100|0489_ , \new_Sorter100|0490_ , \new_Sorter100|0491_ ,
    \new_Sorter100|0492_ , \new_Sorter100|0493_ , \new_Sorter100|0494_ ,
    \new_Sorter100|0495_ , \new_Sorter100|0496_ , \new_Sorter100|0497_ ,
    \new_Sorter100|0498_ , \new_Sorter100|0499_ , \new_Sorter100|0500_ ,
    \new_Sorter100|0599_ , \new_Sorter100|0501_ , \new_Sorter100|0502_ ,
    \new_Sorter100|0503_ , \new_Sorter100|0504_ , \new_Sorter100|0505_ ,
    \new_Sorter100|0506_ , \new_Sorter100|0507_ , \new_Sorter100|0508_ ,
    \new_Sorter100|0509_ , \new_Sorter100|0510_ , \new_Sorter100|0511_ ,
    \new_Sorter100|0512_ , \new_Sorter100|0513_ , \new_Sorter100|0514_ ,
    \new_Sorter100|0515_ , \new_Sorter100|0516_ , \new_Sorter100|0517_ ,
    \new_Sorter100|0518_ , \new_Sorter100|0519_ , \new_Sorter100|0520_ ,
    \new_Sorter100|0521_ , \new_Sorter100|0522_ , \new_Sorter100|0523_ ,
    \new_Sorter100|0524_ , \new_Sorter100|0525_ , \new_Sorter100|0526_ ,
    \new_Sorter100|0527_ , \new_Sorter100|0528_ , \new_Sorter100|0529_ ,
    \new_Sorter100|0530_ , \new_Sorter100|0531_ , \new_Sorter100|0532_ ,
    \new_Sorter100|0533_ , \new_Sorter100|0534_ , \new_Sorter100|0535_ ,
    \new_Sorter100|0536_ , \new_Sorter100|0537_ , \new_Sorter100|0538_ ,
    \new_Sorter100|0539_ , \new_Sorter100|0540_ , \new_Sorter100|0541_ ,
    \new_Sorter100|0542_ , \new_Sorter100|0543_ , \new_Sorter100|0544_ ,
    \new_Sorter100|0545_ , \new_Sorter100|0546_ , \new_Sorter100|0547_ ,
    \new_Sorter100|0548_ , \new_Sorter100|0549_ , \new_Sorter100|0550_ ,
    \new_Sorter100|0551_ , \new_Sorter100|0552_ , \new_Sorter100|0553_ ,
    \new_Sorter100|0554_ , \new_Sorter100|0555_ , \new_Sorter100|0556_ ,
    \new_Sorter100|0557_ , \new_Sorter100|0558_ , \new_Sorter100|0559_ ,
    \new_Sorter100|0560_ , \new_Sorter100|0561_ , \new_Sorter100|0562_ ,
    \new_Sorter100|0563_ , \new_Sorter100|0564_ , \new_Sorter100|0565_ ,
    \new_Sorter100|0566_ , \new_Sorter100|0567_ , \new_Sorter100|0568_ ,
    \new_Sorter100|0569_ , \new_Sorter100|0570_ , \new_Sorter100|0571_ ,
    \new_Sorter100|0572_ , \new_Sorter100|0573_ , \new_Sorter100|0574_ ,
    \new_Sorter100|0575_ , \new_Sorter100|0576_ , \new_Sorter100|0577_ ,
    \new_Sorter100|0578_ , \new_Sorter100|0579_ , \new_Sorter100|0580_ ,
    \new_Sorter100|0581_ , \new_Sorter100|0582_ , \new_Sorter100|0583_ ,
    \new_Sorter100|0584_ , \new_Sorter100|0585_ , \new_Sorter100|0586_ ,
    \new_Sorter100|0587_ , \new_Sorter100|0588_ , \new_Sorter100|0589_ ,
    \new_Sorter100|0590_ , \new_Sorter100|0591_ , \new_Sorter100|0592_ ,
    \new_Sorter100|0593_ , \new_Sorter100|0594_ , \new_Sorter100|0595_ ,
    \new_Sorter100|0596_ , \new_Sorter100|0597_ , \new_Sorter100|0598_ ,
    \new_Sorter100|0600_ , \new_Sorter100|0601_ , \new_Sorter100|0602_ ,
    \new_Sorter100|0603_ , \new_Sorter100|0604_ , \new_Sorter100|0605_ ,
    \new_Sorter100|0606_ , \new_Sorter100|0607_ , \new_Sorter100|0608_ ,
    \new_Sorter100|0609_ , \new_Sorter100|0610_ , \new_Sorter100|0611_ ,
    \new_Sorter100|0612_ , \new_Sorter100|0613_ , \new_Sorter100|0614_ ,
    \new_Sorter100|0615_ , \new_Sorter100|0616_ , \new_Sorter100|0617_ ,
    \new_Sorter100|0618_ , \new_Sorter100|0619_ , \new_Sorter100|0620_ ,
    \new_Sorter100|0621_ , \new_Sorter100|0622_ , \new_Sorter100|0623_ ,
    \new_Sorter100|0624_ , \new_Sorter100|0625_ , \new_Sorter100|0626_ ,
    \new_Sorter100|0627_ , \new_Sorter100|0628_ , \new_Sorter100|0629_ ,
    \new_Sorter100|0630_ , \new_Sorter100|0631_ , \new_Sorter100|0632_ ,
    \new_Sorter100|0633_ , \new_Sorter100|0634_ , \new_Sorter100|0635_ ,
    \new_Sorter100|0636_ , \new_Sorter100|0637_ , \new_Sorter100|0638_ ,
    \new_Sorter100|0639_ , \new_Sorter100|0640_ , \new_Sorter100|0641_ ,
    \new_Sorter100|0642_ , \new_Sorter100|0643_ , \new_Sorter100|0644_ ,
    \new_Sorter100|0645_ , \new_Sorter100|0646_ , \new_Sorter100|0647_ ,
    \new_Sorter100|0648_ , \new_Sorter100|0649_ , \new_Sorter100|0650_ ,
    \new_Sorter100|0651_ , \new_Sorter100|0652_ , \new_Sorter100|0653_ ,
    \new_Sorter100|0654_ , \new_Sorter100|0655_ , \new_Sorter100|0656_ ,
    \new_Sorter100|0657_ , \new_Sorter100|0658_ , \new_Sorter100|0659_ ,
    \new_Sorter100|0660_ , \new_Sorter100|0661_ , \new_Sorter100|0662_ ,
    \new_Sorter100|0663_ , \new_Sorter100|0664_ , \new_Sorter100|0665_ ,
    \new_Sorter100|0666_ , \new_Sorter100|0667_ , \new_Sorter100|0668_ ,
    \new_Sorter100|0669_ , \new_Sorter100|0670_ , \new_Sorter100|0671_ ,
    \new_Sorter100|0672_ , \new_Sorter100|0673_ , \new_Sorter100|0674_ ,
    \new_Sorter100|0675_ , \new_Sorter100|0676_ , \new_Sorter100|0677_ ,
    \new_Sorter100|0678_ , \new_Sorter100|0679_ , \new_Sorter100|0680_ ,
    \new_Sorter100|0681_ , \new_Sorter100|0682_ , \new_Sorter100|0683_ ,
    \new_Sorter100|0684_ , \new_Sorter100|0685_ , \new_Sorter100|0686_ ,
    \new_Sorter100|0687_ , \new_Sorter100|0688_ , \new_Sorter100|0689_ ,
    \new_Sorter100|0690_ , \new_Sorter100|0691_ , \new_Sorter100|0692_ ,
    \new_Sorter100|0693_ , \new_Sorter100|0694_ , \new_Sorter100|0695_ ,
    \new_Sorter100|0696_ , \new_Sorter100|0697_ , \new_Sorter100|0698_ ,
    \new_Sorter100|0699_ , \new_Sorter100|0700_ , \new_Sorter100|0799_ ,
    \new_Sorter100|0701_ , \new_Sorter100|0702_ , \new_Sorter100|0703_ ,
    \new_Sorter100|0704_ , \new_Sorter100|0705_ , \new_Sorter100|0706_ ,
    \new_Sorter100|0707_ , \new_Sorter100|0708_ , \new_Sorter100|0709_ ,
    \new_Sorter100|0710_ , \new_Sorter100|0711_ , \new_Sorter100|0712_ ,
    \new_Sorter100|0713_ , \new_Sorter100|0714_ , \new_Sorter100|0715_ ,
    \new_Sorter100|0716_ , \new_Sorter100|0717_ , \new_Sorter100|0718_ ,
    \new_Sorter100|0719_ , \new_Sorter100|0720_ , \new_Sorter100|0721_ ,
    \new_Sorter100|0722_ , \new_Sorter100|0723_ , \new_Sorter100|0724_ ,
    \new_Sorter100|0725_ , \new_Sorter100|0726_ , \new_Sorter100|0727_ ,
    \new_Sorter100|0728_ , \new_Sorter100|0729_ , \new_Sorter100|0730_ ,
    \new_Sorter100|0731_ , \new_Sorter100|0732_ , \new_Sorter100|0733_ ,
    \new_Sorter100|0734_ , \new_Sorter100|0735_ , \new_Sorter100|0736_ ,
    \new_Sorter100|0737_ , \new_Sorter100|0738_ , \new_Sorter100|0739_ ,
    \new_Sorter100|0740_ , \new_Sorter100|0741_ , \new_Sorter100|0742_ ,
    \new_Sorter100|0743_ , \new_Sorter100|0744_ , \new_Sorter100|0745_ ,
    \new_Sorter100|0746_ , \new_Sorter100|0747_ , \new_Sorter100|0748_ ,
    \new_Sorter100|0749_ , \new_Sorter100|0750_ , \new_Sorter100|0751_ ,
    \new_Sorter100|0752_ , \new_Sorter100|0753_ , \new_Sorter100|0754_ ,
    \new_Sorter100|0755_ , \new_Sorter100|0756_ , \new_Sorter100|0757_ ,
    \new_Sorter100|0758_ , \new_Sorter100|0759_ , \new_Sorter100|0760_ ,
    \new_Sorter100|0761_ , \new_Sorter100|0762_ , \new_Sorter100|0763_ ,
    \new_Sorter100|0764_ , \new_Sorter100|0765_ , \new_Sorter100|0766_ ,
    \new_Sorter100|0767_ , \new_Sorter100|0768_ , \new_Sorter100|0769_ ,
    \new_Sorter100|0770_ , \new_Sorter100|0771_ , \new_Sorter100|0772_ ,
    \new_Sorter100|0773_ , \new_Sorter100|0774_ , \new_Sorter100|0775_ ,
    \new_Sorter100|0776_ , \new_Sorter100|0777_ , \new_Sorter100|0778_ ,
    \new_Sorter100|0779_ , \new_Sorter100|0780_ , \new_Sorter100|0781_ ,
    \new_Sorter100|0782_ , \new_Sorter100|0783_ , \new_Sorter100|0784_ ,
    \new_Sorter100|0785_ , \new_Sorter100|0786_ , \new_Sorter100|0787_ ,
    \new_Sorter100|0788_ , \new_Sorter100|0789_ , \new_Sorter100|0790_ ,
    \new_Sorter100|0791_ , \new_Sorter100|0792_ , \new_Sorter100|0793_ ,
    \new_Sorter100|0794_ , \new_Sorter100|0795_ , \new_Sorter100|0796_ ,
    \new_Sorter100|0797_ , \new_Sorter100|0798_ , \new_Sorter100|0800_ ,
    \new_Sorter100|0801_ , \new_Sorter100|0802_ , \new_Sorter100|0803_ ,
    \new_Sorter100|0804_ , \new_Sorter100|0805_ , \new_Sorter100|0806_ ,
    \new_Sorter100|0807_ , \new_Sorter100|0808_ , \new_Sorter100|0809_ ,
    \new_Sorter100|0810_ , \new_Sorter100|0811_ , \new_Sorter100|0812_ ,
    \new_Sorter100|0813_ , \new_Sorter100|0814_ , \new_Sorter100|0815_ ,
    \new_Sorter100|0816_ , \new_Sorter100|0817_ , \new_Sorter100|0818_ ,
    \new_Sorter100|0819_ , \new_Sorter100|0820_ , \new_Sorter100|0821_ ,
    \new_Sorter100|0822_ , \new_Sorter100|0823_ , \new_Sorter100|0824_ ,
    \new_Sorter100|0825_ , \new_Sorter100|0826_ , \new_Sorter100|0827_ ,
    \new_Sorter100|0828_ , \new_Sorter100|0829_ , \new_Sorter100|0830_ ,
    \new_Sorter100|0831_ , \new_Sorter100|0832_ , \new_Sorter100|0833_ ,
    \new_Sorter100|0834_ , \new_Sorter100|0835_ , \new_Sorter100|0836_ ,
    \new_Sorter100|0837_ , \new_Sorter100|0838_ , \new_Sorter100|0839_ ,
    \new_Sorter100|0840_ , \new_Sorter100|0841_ , \new_Sorter100|0842_ ,
    \new_Sorter100|0843_ , \new_Sorter100|0844_ , \new_Sorter100|0845_ ,
    \new_Sorter100|0846_ , \new_Sorter100|0847_ , \new_Sorter100|0848_ ,
    \new_Sorter100|0849_ , \new_Sorter100|0850_ , \new_Sorter100|0851_ ,
    \new_Sorter100|0852_ , \new_Sorter100|0853_ , \new_Sorter100|0854_ ,
    \new_Sorter100|0855_ , \new_Sorter100|0856_ , \new_Sorter100|0857_ ,
    \new_Sorter100|0858_ , \new_Sorter100|0859_ , \new_Sorter100|0860_ ,
    \new_Sorter100|0861_ , \new_Sorter100|0862_ , \new_Sorter100|0863_ ,
    \new_Sorter100|0864_ , \new_Sorter100|0865_ , \new_Sorter100|0866_ ,
    \new_Sorter100|0867_ , \new_Sorter100|0868_ , \new_Sorter100|0869_ ,
    \new_Sorter100|0870_ , \new_Sorter100|0871_ , \new_Sorter100|0872_ ,
    \new_Sorter100|0873_ , \new_Sorter100|0874_ , \new_Sorter100|0875_ ,
    \new_Sorter100|0876_ , \new_Sorter100|0877_ , \new_Sorter100|0878_ ,
    \new_Sorter100|0879_ , \new_Sorter100|0880_ , \new_Sorter100|0881_ ,
    \new_Sorter100|0882_ , \new_Sorter100|0883_ , \new_Sorter100|0884_ ,
    \new_Sorter100|0885_ , \new_Sorter100|0886_ , \new_Sorter100|0887_ ,
    \new_Sorter100|0888_ , \new_Sorter100|0889_ , \new_Sorter100|0890_ ,
    \new_Sorter100|0891_ , \new_Sorter100|0892_ , \new_Sorter100|0893_ ,
    \new_Sorter100|0894_ , \new_Sorter100|0895_ , \new_Sorter100|0896_ ,
    \new_Sorter100|0897_ , \new_Sorter100|0898_ , \new_Sorter100|0899_ ,
    \new_Sorter100|0900_ , \new_Sorter100|0999_ , \new_Sorter100|0901_ ,
    \new_Sorter100|0902_ , \new_Sorter100|0903_ , \new_Sorter100|0904_ ,
    \new_Sorter100|0905_ , \new_Sorter100|0906_ , \new_Sorter100|0907_ ,
    \new_Sorter100|0908_ , \new_Sorter100|0909_ , \new_Sorter100|0910_ ,
    \new_Sorter100|0911_ , \new_Sorter100|0912_ , \new_Sorter100|0913_ ,
    \new_Sorter100|0914_ , \new_Sorter100|0915_ , \new_Sorter100|0916_ ,
    \new_Sorter100|0917_ , \new_Sorter100|0918_ , \new_Sorter100|0919_ ,
    \new_Sorter100|0920_ , \new_Sorter100|0921_ , \new_Sorter100|0922_ ,
    \new_Sorter100|0923_ , \new_Sorter100|0924_ , \new_Sorter100|0925_ ,
    \new_Sorter100|0926_ , \new_Sorter100|0927_ , \new_Sorter100|0928_ ,
    \new_Sorter100|0929_ , \new_Sorter100|0930_ , \new_Sorter100|0931_ ,
    \new_Sorter100|0932_ , \new_Sorter100|0933_ , \new_Sorter100|0934_ ,
    \new_Sorter100|0935_ , \new_Sorter100|0936_ , \new_Sorter100|0937_ ,
    \new_Sorter100|0938_ , \new_Sorter100|0939_ , \new_Sorter100|0940_ ,
    \new_Sorter100|0941_ , \new_Sorter100|0942_ , \new_Sorter100|0943_ ,
    \new_Sorter100|0944_ , \new_Sorter100|0945_ , \new_Sorter100|0946_ ,
    \new_Sorter100|0947_ , \new_Sorter100|0948_ , \new_Sorter100|0949_ ,
    \new_Sorter100|0950_ , \new_Sorter100|0951_ , \new_Sorter100|0952_ ,
    \new_Sorter100|0953_ , \new_Sorter100|0954_ , \new_Sorter100|0955_ ,
    \new_Sorter100|0956_ , \new_Sorter100|0957_ , \new_Sorter100|0958_ ,
    \new_Sorter100|0959_ , \new_Sorter100|0960_ , \new_Sorter100|0961_ ,
    \new_Sorter100|0962_ , \new_Sorter100|0963_ , \new_Sorter100|0964_ ,
    \new_Sorter100|0965_ , \new_Sorter100|0966_ , \new_Sorter100|0967_ ,
    \new_Sorter100|0968_ , \new_Sorter100|0969_ , \new_Sorter100|0970_ ,
    \new_Sorter100|0971_ , \new_Sorter100|0972_ , \new_Sorter100|0973_ ,
    \new_Sorter100|0974_ , \new_Sorter100|0975_ , \new_Sorter100|0976_ ,
    \new_Sorter100|0977_ , \new_Sorter100|0978_ , \new_Sorter100|0979_ ,
    \new_Sorter100|0980_ , \new_Sorter100|0981_ , \new_Sorter100|0982_ ,
    \new_Sorter100|0983_ , \new_Sorter100|0984_ , \new_Sorter100|0985_ ,
    \new_Sorter100|0986_ , \new_Sorter100|0987_ , \new_Sorter100|0988_ ,
    \new_Sorter100|0989_ , \new_Sorter100|0990_ , \new_Sorter100|0991_ ,
    \new_Sorter100|0992_ , \new_Sorter100|0993_ , \new_Sorter100|0994_ ,
    \new_Sorter100|0995_ , \new_Sorter100|0996_ , \new_Sorter100|0997_ ,
    \new_Sorter100|0998_ , \new_Sorter100|1000_ , \new_Sorter100|1001_ ,
    \new_Sorter100|1002_ , \new_Sorter100|1003_ , \new_Sorter100|1004_ ,
    \new_Sorter100|1005_ , \new_Sorter100|1006_ , \new_Sorter100|1007_ ,
    \new_Sorter100|1008_ , \new_Sorter100|1009_ , \new_Sorter100|1010_ ,
    \new_Sorter100|1011_ , \new_Sorter100|1012_ , \new_Sorter100|1013_ ,
    \new_Sorter100|1014_ , \new_Sorter100|1015_ , \new_Sorter100|1016_ ,
    \new_Sorter100|1017_ , \new_Sorter100|1018_ , \new_Sorter100|1019_ ,
    \new_Sorter100|1020_ , \new_Sorter100|1021_ , \new_Sorter100|1022_ ,
    \new_Sorter100|1023_ , \new_Sorter100|1024_ , \new_Sorter100|1025_ ,
    \new_Sorter100|1026_ , \new_Sorter100|1027_ , \new_Sorter100|1028_ ,
    \new_Sorter100|1029_ , \new_Sorter100|1030_ , \new_Sorter100|1031_ ,
    \new_Sorter100|1032_ , \new_Sorter100|1033_ , \new_Sorter100|1034_ ,
    \new_Sorter100|1035_ , \new_Sorter100|1036_ , \new_Sorter100|1037_ ,
    \new_Sorter100|1038_ , \new_Sorter100|1039_ , \new_Sorter100|1040_ ,
    \new_Sorter100|1041_ , \new_Sorter100|1042_ , \new_Sorter100|1043_ ,
    \new_Sorter100|1044_ , \new_Sorter100|1045_ , \new_Sorter100|1046_ ,
    \new_Sorter100|1047_ , \new_Sorter100|1048_ , \new_Sorter100|1049_ ,
    \new_Sorter100|1050_ , \new_Sorter100|1051_ , \new_Sorter100|1052_ ,
    \new_Sorter100|1053_ , \new_Sorter100|1054_ , \new_Sorter100|1055_ ,
    \new_Sorter100|1056_ , \new_Sorter100|1057_ , \new_Sorter100|1058_ ,
    \new_Sorter100|1059_ , \new_Sorter100|1060_ , \new_Sorter100|1061_ ,
    \new_Sorter100|1062_ , \new_Sorter100|1063_ , \new_Sorter100|1064_ ,
    \new_Sorter100|1065_ , \new_Sorter100|1066_ , \new_Sorter100|1067_ ,
    \new_Sorter100|1068_ , \new_Sorter100|1069_ , \new_Sorter100|1070_ ,
    \new_Sorter100|1071_ , \new_Sorter100|1072_ , \new_Sorter100|1073_ ,
    \new_Sorter100|1074_ , \new_Sorter100|1075_ , \new_Sorter100|1076_ ,
    \new_Sorter100|1077_ , \new_Sorter100|1078_ , \new_Sorter100|1079_ ,
    \new_Sorter100|1080_ , \new_Sorter100|1081_ , \new_Sorter100|1082_ ,
    \new_Sorter100|1083_ , \new_Sorter100|1084_ , \new_Sorter100|1085_ ,
    \new_Sorter100|1086_ , \new_Sorter100|1087_ , \new_Sorter100|1088_ ,
    \new_Sorter100|1089_ , \new_Sorter100|1090_ , \new_Sorter100|1091_ ,
    \new_Sorter100|1092_ , \new_Sorter100|1093_ , \new_Sorter100|1094_ ,
    \new_Sorter100|1095_ , \new_Sorter100|1096_ , \new_Sorter100|1097_ ,
    \new_Sorter100|1098_ , \new_Sorter100|1099_ , \new_Sorter100|1100_ ,
    \new_Sorter100|1199_ , \new_Sorter100|1101_ , \new_Sorter100|1102_ ,
    \new_Sorter100|1103_ , \new_Sorter100|1104_ , \new_Sorter100|1105_ ,
    \new_Sorter100|1106_ , \new_Sorter100|1107_ , \new_Sorter100|1108_ ,
    \new_Sorter100|1109_ , \new_Sorter100|1110_ , \new_Sorter100|1111_ ,
    \new_Sorter100|1112_ , \new_Sorter100|1113_ , \new_Sorter100|1114_ ,
    \new_Sorter100|1115_ , \new_Sorter100|1116_ , \new_Sorter100|1117_ ,
    \new_Sorter100|1118_ , \new_Sorter100|1119_ , \new_Sorter100|1120_ ,
    \new_Sorter100|1121_ , \new_Sorter100|1122_ , \new_Sorter100|1123_ ,
    \new_Sorter100|1124_ , \new_Sorter100|1125_ , \new_Sorter100|1126_ ,
    \new_Sorter100|1127_ , \new_Sorter100|1128_ , \new_Sorter100|1129_ ,
    \new_Sorter100|1130_ , \new_Sorter100|1131_ , \new_Sorter100|1132_ ,
    \new_Sorter100|1133_ , \new_Sorter100|1134_ , \new_Sorter100|1135_ ,
    \new_Sorter100|1136_ , \new_Sorter100|1137_ , \new_Sorter100|1138_ ,
    \new_Sorter100|1139_ , \new_Sorter100|1140_ , \new_Sorter100|1141_ ,
    \new_Sorter100|1142_ , \new_Sorter100|1143_ , \new_Sorter100|1144_ ,
    \new_Sorter100|1145_ , \new_Sorter100|1146_ , \new_Sorter100|1147_ ,
    \new_Sorter100|1148_ , \new_Sorter100|1149_ , \new_Sorter100|1150_ ,
    \new_Sorter100|1151_ , \new_Sorter100|1152_ , \new_Sorter100|1153_ ,
    \new_Sorter100|1154_ , \new_Sorter100|1155_ , \new_Sorter100|1156_ ,
    \new_Sorter100|1157_ , \new_Sorter100|1158_ , \new_Sorter100|1159_ ,
    \new_Sorter100|1160_ , \new_Sorter100|1161_ , \new_Sorter100|1162_ ,
    \new_Sorter100|1163_ , \new_Sorter100|1164_ , \new_Sorter100|1165_ ,
    \new_Sorter100|1166_ , \new_Sorter100|1167_ , \new_Sorter100|1168_ ,
    \new_Sorter100|1169_ , \new_Sorter100|1170_ , \new_Sorter100|1171_ ,
    \new_Sorter100|1172_ , \new_Sorter100|1173_ , \new_Sorter100|1174_ ,
    \new_Sorter100|1175_ , \new_Sorter100|1176_ , \new_Sorter100|1177_ ,
    \new_Sorter100|1178_ , \new_Sorter100|1179_ , \new_Sorter100|1180_ ,
    \new_Sorter100|1181_ , \new_Sorter100|1182_ , \new_Sorter100|1183_ ,
    \new_Sorter100|1184_ , \new_Sorter100|1185_ , \new_Sorter100|1186_ ,
    \new_Sorter100|1187_ , \new_Sorter100|1188_ , \new_Sorter100|1189_ ,
    \new_Sorter100|1190_ , \new_Sorter100|1191_ , \new_Sorter100|1192_ ,
    \new_Sorter100|1193_ , \new_Sorter100|1194_ , \new_Sorter100|1195_ ,
    \new_Sorter100|1196_ , \new_Sorter100|1197_ , \new_Sorter100|1198_ ,
    \new_Sorter100|1200_ , \new_Sorter100|1201_ , \new_Sorter100|1202_ ,
    \new_Sorter100|1203_ , \new_Sorter100|1204_ , \new_Sorter100|1205_ ,
    \new_Sorter100|1206_ , \new_Sorter100|1207_ , \new_Sorter100|1208_ ,
    \new_Sorter100|1209_ , \new_Sorter100|1210_ , \new_Sorter100|1211_ ,
    \new_Sorter100|1212_ , \new_Sorter100|1213_ , \new_Sorter100|1214_ ,
    \new_Sorter100|1215_ , \new_Sorter100|1216_ , \new_Sorter100|1217_ ,
    \new_Sorter100|1218_ , \new_Sorter100|1219_ , \new_Sorter100|1220_ ,
    \new_Sorter100|1221_ , \new_Sorter100|1222_ , \new_Sorter100|1223_ ,
    \new_Sorter100|1224_ , \new_Sorter100|1225_ , \new_Sorter100|1226_ ,
    \new_Sorter100|1227_ , \new_Sorter100|1228_ , \new_Sorter100|1229_ ,
    \new_Sorter100|1230_ , \new_Sorter100|1231_ , \new_Sorter100|1232_ ,
    \new_Sorter100|1233_ , \new_Sorter100|1234_ , \new_Sorter100|1235_ ,
    \new_Sorter100|1236_ , \new_Sorter100|1237_ , \new_Sorter100|1238_ ,
    \new_Sorter100|1239_ , \new_Sorter100|1240_ , \new_Sorter100|1241_ ,
    \new_Sorter100|1242_ , \new_Sorter100|1243_ , \new_Sorter100|1244_ ,
    \new_Sorter100|1245_ , \new_Sorter100|1246_ , \new_Sorter100|1247_ ,
    \new_Sorter100|1248_ , \new_Sorter100|1249_ , \new_Sorter100|1250_ ,
    \new_Sorter100|1251_ , \new_Sorter100|1252_ , \new_Sorter100|1253_ ,
    \new_Sorter100|1254_ , \new_Sorter100|1255_ , \new_Sorter100|1256_ ,
    \new_Sorter100|1257_ , \new_Sorter100|1258_ , \new_Sorter100|1259_ ,
    \new_Sorter100|1260_ , \new_Sorter100|1261_ , \new_Sorter100|1262_ ,
    \new_Sorter100|1263_ , \new_Sorter100|1264_ , \new_Sorter100|1265_ ,
    \new_Sorter100|1266_ , \new_Sorter100|1267_ , \new_Sorter100|1268_ ,
    \new_Sorter100|1269_ , \new_Sorter100|1270_ , \new_Sorter100|1271_ ,
    \new_Sorter100|1272_ , \new_Sorter100|1273_ , \new_Sorter100|1274_ ,
    \new_Sorter100|1275_ , \new_Sorter100|1276_ , \new_Sorter100|1277_ ,
    \new_Sorter100|1278_ , \new_Sorter100|1279_ , \new_Sorter100|1280_ ,
    \new_Sorter100|1281_ , \new_Sorter100|1282_ , \new_Sorter100|1283_ ,
    \new_Sorter100|1284_ , \new_Sorter100|1285_ , \new_Sorter100|1286_ ,
    \new_Sorter100|1287_ , \new_Sorter100|1288_ , \new_Sorter100|1289_ ,
    \new_Sorter100|1290_ , \new_Sorter100|1291_ , \new_Sorter100|1292_ ,
    \new_Sorter100|1293_ , \new_Sorter100|1294_ , \new_Sorter100|1295_ ,
    \new_Sorter100|1296_ , \new_Sorter100|1297_ , \new_Sorter100|1298_ ,
    \new_Sorter100|1299_ , \new_Sorter100|1300_ , \new_Sorter100|1399_ ,
    \new_Sorter100|1301_ , \new_Sorter100|1302_ , \new_Sorter100|1303_ ,
    \new_Sorter100|1304_ , \new_Sorter100|1305_ , \new_Sorter100|1306_ ,
    \new_Sorter100|1307_ , \new_Sorter100|1308_ , \new_Sorter100|1309_ ,
    \new_Sorter100|1310_ , \new_Sorter100|1311_ , \new_Sorter100|1312_ ,
    \new_Sorter100|1313_ , \new_Sorter100|1314_ , \new_Sorter100|1315_ ,
    \new_Sorter100|1316_ , \new_Sorter100|1317_ , \new_Sorter100|1318_ ,
    \new_Sorter100|1319_ , \new_Sorter100|1320_ , \new_Sorter100|1321_ ,
    \new_Sorter100|1322_ , \new_Sorter100|1323_ , \new_Sorter100|1324_ ,
    \new_Sorter100|1325_ , \new_Sorter100|1326_ , \new_Sorter100|1327_ ,
    \new_Sorter100|1328_ , \new_Sorter100|1329_ , \new_Sorter100|1330_ ,
    \new_Sorter100|1331_ , \new_Sorter100|1332_ , \new_Sorter100|1333_ ,
    \new_Sorter100|1334_ , \new_Sorter100|1335_ , \new_Sorter100|1336_ ,
    \new_Sorter100|1337_ , \new_Sorter100|1338_ , \new_Sorter100|1339_ ,
    \new_Sorter100|1340_ , \new_Sorter100|1341_ , \new_Sorter100|1342_ ,
    \new_Sorter100|1343_ , \new_Sorter100|1344_ , \new_Sorter100|1345_ ,
    \new_Sorter100|1346_ , \new_Sorter100|1347_ , \new_Sorter100|1348_ ,
    \new_Sorter100|1349_ , \new_Sorter100|1350_ , \new_Sorter100|1351_ ,
    \new_Sorter100|1352_ , \new_Sorter100|1353_ , \new_Sorter100|1354_ ,
    \new_Sorter100|1355_ , \new_Sorter100|1356_ , \new_Sorter100|1357_ ,
    \new_Sorter100|1358_ , \new_Sorter100|1359_ , \new_Sorter100|1360_ ,
    \new_Sorter100|1361_ , \new_Sorter100|1362_ , \new_Sorter100|1363_ ,
    \new_Sorter100|1364_ , \new_Sorter100|1365_ , \new_Sorter100|1366_ ,
    \new_Sorter100|1367_ , \new_Sorter100|1368_ , \new_Sorter100|1369_ ,
    \new_Sorter100|1370_ , \new_Sorter100|1371_ , \new_Sorter100|1372_ ,
    \new_Sorter100|1373_ , \new_Sorter100|1374_ , \new_Sorter100|1375_ ,
    \new_Sorter100|1376_ , \new_Sorter100|1377_ , \new_Sorter100|1378_ ,
    \new_Sorter100|1379_ , \new_Sorter100|1380_ , \new_Sorter100|1381_ ,
    \new_Sorter100|1382_ , \new_Sorter100|1383_ , \new_Sorter100|1384_ ,
    \new_Sorter100|1385_ , \new_Sorter100|1386_ , \new_Sorter100|1387_ ,
    \new_Sorter100|1388_ , \new_Sorter100|1389_ , \new_Sorter100|1390_ ,
    \new_Sorter100|1391_ , \new_Sorter100|1392_ , \new_Sorter100|1393_ ,
    \new_Sorter100|1394_ , \new_Sorter100|1395_ , \new_Sorter100|1396_ ,
    \new_Sorter100|1397_ , \new_Sorter100|1398_ , \new_Sorter100|1400_ ,
    \new_Sorter100|1401_ , \new_Sorter100|1402_ , \new_Sorter100|1403_ ,
    \new_Sorter100|1404_ , \new_Sorter100|1405_ , \new_Sorter100|1406_ ,
    \new_Sorter100|1407_ , \new_Sorter100|1408_ , \new_Sorter100|1409_ ,
    \new_Sorter100|1410_ , \new_Sorter100|1411_ , \new_Sorter100|1412_ ,
    \new_Sorter100|1413_ , \new_Sorter100|1414_ , \new_Sorter100|1415_ ,
    \new_Sorter100|1416_ , \new_Sorter100|1417_ , \new_Sorter100|1418_ ,
    \new_Sorter100|1419_ , \new_Sorter100|1420_ , \new_Sorter100|1421_ ,
    \new_Sorter100|1422_ , \new_Sorter100|1423_ , \new_Sorter100|1424_ ,
    \new_Sorter100|1425_ , \new_Sorter100|1426_ , \new_Sorter100|1427_ ,
    \new_Sorter100|1428_ , \new_Sorter100|1429_ , \new_Sorter100|1430_ ,
    \new_Sorter100|1431_ , \new_Sorter100|1432_ , \new_Sorter100|1433_ ,
    \new_Sorter100|1434_ , \new_Sorter100|1435_ , \new_Sorter100|1436_ ,
    \new_Sorter100|1437_ , \new_Sorter100|1438_ , \new_Sorter100|1439_ ,
    \new_Sorter100|1440_ , \new_Sorter100|1441_ , \new_Sorter100|1442_ ,
    \new_Sorter100|1443_ , \new_Sorter100|1444_ , \new_Sorter100|1445_ ,
    \new_Sorter100|1446_ , \new_Sorter100|1447_ , \new_Sorter100|1448_ ,
    \new_Sorter100|1449_ , \new_Sorter100|1450_ , \new_Sorter100|1451_ ,
    \new_Sorter100|1452_ , \new_Sorter100|1453_ , \new_Sorter100|1454_ ,
    \new_Sorter100|1455_ , \new_Sorter100|1456_ , \new_Sorter100|1457_ ,
    \new_Sorter100|1458_ , \new_Sorter100|1459_ , \new_Sorter100|1460_ ,
    \new_Sorter100|1461_ , \new_Sorter100|1462_ , \new_Sorter100|1463_ ,
    \new_Sorter100|1464_ , \new_Sorter100|1465_ , \new_Sorter100|1466_ ,
    \new_Sorter100|1467_ , \new_Sorter100|1468_ , \new_Sorter100|1469_ ,
    \new_Sorter100|1470_ , \new_Sorter100|1471_ , \new_Sorter100|1472_ ,
    \new_Sorter100|1473_ , \new_Sorter100|1474_ , \new_Sorter100|1475_ ,
    \new_Sorter100|1476_ , \new_Sorter100|1477_ , \new_Sorter100|1478_ ,
    \new_Sorter100|1479_ , \new_Sorter100|1480_ , \new_Sorter100|1481_ ,
    \new_Sorter100|1482_ , \new_Sorter100|1483_ , \new_Sorter100|1484_ ,
    \new_Sorter100|1485_ , \new_Sorter100|1486_ , \new_Sorter100|1487_ ,
    \new_Sorter100|1488_ , \new_Sorter100|1489_ , \new_Sorter100|1490_ ,
    \new_Sorter100|1491_ , \new_Sorter100|1492_ , \new_Sorter100|1493_ ,
    \new_Sorter100|1494_ , \new_Sorter100|1495_ , \new_Sorter100|1496_ ,
    \new_Sorter100|1497_ , \new_Sorter100|1498_ , \new_Sorter100|1499_ ,
    \new_Sorter100|1500_ , \new_Sorter100|1599_ , \new_Sorter100|1501_ ,
    \new_Sorter100|1502_ , \new_Sorter100|1503_ , \new_Sorter100|1504_ ,
    \new_Sorter100|1505_ , \new_Sorter100|1506_ , \new_Sorter100|1507_ ,
    \new_Sorter100|1508_ , \new_Sorter100|1509_ , \new_Sorter100|1510_ ,
    \new_Sorter100|1511_ , \new_Sorter100|1512_ , \new_Sorter100|1513_ ,
    \new_Sorter100|1514_ , \new_Sorter100|1515_ , \new_Sorter100|1516_ ,
    \new_Sorter100|1517_ , \new_Sorter100|1518_ , \new_Sorter100|1519_ ,
    \new_Sorter100|1520_ , \new_Sorter100|1521_ , \new_Sorter100|1522_ ,
    \new_Sorter100|1523_ , \new_Sorter100|1524_ , \new_Sorter100|1525_ ,
    \new_Sorter100|1526_ , \new_Sorter100|1527_ , \new_Sorter100|1528_ ,
    \new_Sorter100|1529_ , \new_Sorter100|1530_ , \new_Sorter100|1531_ ,
    \new_Sorter100|1532_ , \new_Sorter100|1533_ , \new_Sorter100|1534_ ,
    \new_Sorter100|1535_ , \new_Sorter100|1536_ , \new_Sorter100|1537_ ,
    \new_Sorter100|1538_ , \new_Sorter100|1539_ , \new_Sorter100|1540_ ,
    \new_Sorter100|1541_ , \new_Sorter100|1542_ , \new_Sorter100|1543_ ,
    \new_Sorter100|1544_ , \new_Sorter100|1545_ , \new_Sorter100|1546_ ,
    \new_Sorter100|1547_ , \new_Sorter100|1548_ , \new_Sorter100|1549_ ,
    \new_Sorter100|1550_ , \new_Sorter100|1551_ , \new_Sorter100|1552_ ,
    \new_Sorter100|1553_ , \new_Sorter100|1554_ , \new_Sorter100|1555_ ,
    \new_Sorter100|1556_ , \new_Sorter100|1557_ , \new_Sorter100|1558_ ,
    \new_Sorter100|1559_ , \new_Sorter100|1560_ , \new_Sorter100|1561_ ,
    \new_Sorter100|1562_ , \new_Sorter100|1563_ , \new_Sorter100|1564_ ,
    \new_Sorter100|1565_ , \new_Sorter100|1566_ , \new_Sorter100|1567_ ,
    \new_Sorter100|1568_ , \new_Sorter100|1569_ , \new_Sorter100|1570_ ,
    \new_Sorter100|1571_ , \new_Sorter100|1572_ , \new_Sorter100|1573_ ,
    \new_Sorter100|1574_ , \new_Sorter100|1575_ , \new_Sorter100|1576_ ,
    \new_Sorter100|1577_ , \new_Sorter100|1578_ , \new_Sorter100|1579_ ,
    \new_Sorter100|1580_ , \new_Sorter100|1581_ , \new_Sorter100|1582_ ,
    \new_Sorter100|1583_ , \new_Sorter100|1584_ , \new_Sorter100|1585_ ,
    \new_Sorter100|1586_ , \new_Sorter100|1587_ , \new_Sorter100|1588_ ,
    \new_Sorter100|1589_ , \new_Sorter100|1590_ , \new_Sorter100|1591_ ,
    \new_Sorter100|1592_ , \new_Sorter100|1593_ , \new_Sorter100|1594_ ,
    \new_Sorter100|1595_ , \new_Sorter100|1596_ , \new_Sorter100|1597_ ,
    \new_Sorter100|1598_ , \new_Sorter100|1600_ , \new_Sorter100|1601_ ,
    \new_Sorter100|1602_ , \new_Sorter100|1603_ , \new_Sorter100|1604_ ,
    \new_Sorter100|1605_ , \new_Sorter100|1606_ , \new_Sorter100|1607_ ,
    \new_Sorter100|1608_ , \new_Sorter100|1609_ , \new_Sorter100|1610_ ,
    \new_Sorter100|1611_ , \new_Sorter100|1612_ , \new_Sorter100|1613_ ,
    \new_Sorter100|1614_ , \new_Sorter100|1615_ , \new_Sorter100|1616_ ,
    \new_Sorter100|1617_ , \new_Sorter100|1618_ , \new_Sorter100|1619_ ,
    \new_Sorter100|1620_ , \new_Sorter100|1621_ , \new_Sorter100|1622_ ,
    \new_Sorter100|1623_ , \new_Sorter100|1624_ , \new_Sorter100|1625_ ,
    \new_Sorter100|1626_ , \new_Sorter100|1627_ , \new_Sorter100|1628_ ,
    \new_Sorter100|1629_ , \new_Sorter100|1630_ , \new_Sorter100|1631_ ,
    \new_Sorter100|1632_ , \new_Sorter100|1633_ , \new_Sorter100|1634_ ,
    \new_Sorter100|1635_ , \new_Sorter100|1636_ , \new_Sorter100|1637_ ,
    \new_Sorter100|1638_ , \new_Sorter100|1639_ , \new_Sorter100|1640_ ,
    \new_Sorter100|1641_ , \new_Sorter100|1642_ , \new_Sorter100|1643_ ,
    \new_Sorter100|1644_ , \new_Sorter100|1645_ , \new_Sorter100|1646_ ,
    \new_Sorter100|1647_ , \new_Sorter100|1648_ , \new_Sorter100|1649_ ,
    \new_Sorter100|1650_ , \new_Sorter100|1651_ , \new_Sorter100|1652_ ,
    \new_Sorter100|1653_ , \new_Sorter100|1654_ , \new_Sorter100|1655_ ,
    \new_Sorter100|1656_ , \new_Sorter100|1657_ , \new_Sorter100|1658_ ,
    \new_Sorter100|1659_ , \new_Sorter100|1660_ , \new_Sorter100|1661_ ,
    \new_Sorter100|1662_ , \new_Sorter100|1663_ , \new_Sorter100|1664_ ,
    \new_Sorter100|1665_ , \new_Sorter100|1666_ , \new_Sorter100|1667_ ,
    \new_Sorter100|1668_ , \new_Sorter100|1669_ , \new_Sorter100|1670_ ,
    \new_Sorter100|1671_ , \new_Sorter100|1672_ , \new_Sorter100|1673_ ,
    \new_Sorter100|1674_ , \new_Sorter100|1675_ , \new_Sorter100|1676_ ,
    \new_Sorter100|1677_ , \new_Sorter100|1678_ , \new_Sorter100|1679_ ,
    \new_Sorter100|1680_ , \new_Sorter100|1681_ , \new_Sorter100|1682_ ,
    \new_Sorter100|1683_ , \new_Sorter100|1684_ , \new_Sorter100|1685_ ,
    \new_Sorter100|1686_ , \new_Sorter100|1687_ , \new_Sorter100|1688_ ,
    \new_Sorter100|1689_ , \new_Sorter100|1690_ , \new_Sorter100|1691_ ,
    \new_Sorter100|1692_ , \new_Sorter100|1693_ , \new_Sorter100|1694_ ,
    \new_Sorter100|1695_ , \new_Sorter100|1696_ , \new_Sorter100|1697_ ,
    \new_Sorter100|1698_ , \new_Sorter100|1699_ , \new_Sorter100|1700_ ,
    \new_Sorter100|1799_ , \new_Sorter100|1701_ , \new_Sorter100|1702_ ,
    \new_Sorter100|1703_ , \new_Sorter100|1704_ , \new_Sorter100|1705_ ,
    \new_Sorter100|1706_ , \new_Sorter100|1707_ , \new_Sorter100|1708_ ,
    \new_Sorter100|1709_ , \new_Sorter100|1710_ , \new_Sorter100|1711_ ,
    \new_Sorter100|1712_ , \new_Sorter100|1713_ , \new_Sorter100|1714_ ,
    \new_Sorter100|1715_ , \new_Sorter100|1716_ , \new_Sorter100|1717_ ,
    \new_Sorter100|1718_ , \new_Sorter100|1719_ , \new_Sorter100|1720_ ,
    \new_Sorter100|1721_ , \new_Sorter100|1722_ , \new_Sorter100|1723_ ,
    \new_Sorter100|1724_ , \new_Sorter100|1725_ , \new_Sorter100|1726_ ,
    \new_Sorter100|1727_ , \new_Sorter100|1728_ , \new_Sorter100|1729_ ,
    \new_Sorter100|1730_ , \new_Sorter100|1731_ , \new_Sorter100|1732_ ,
    \new_Sorter100|1733_ , \new_Sorter100|1734_ , \new_Sorter100|1735_ ,
    \new_Sorter100|1736_ , \new_Sorter100|1737_ , \new_Sorter100|1738_ ,
    \new_Sorter100|1739_ , \new_Sorter100|1740_ , \new_Sorter100|1741_ ,
    \new_Sorter100|1742_ , \new_Sorter100|1743_ , \new_Sorter100|1744_ ,
    \new_Sorter100|1745_ , \new_Sorter100|1746_ , \new_Sorter100|1747_ ,
    \new_Sorter100|1748_ , \new_Sorter100|1749_ , \new_Sorter100|1750_ ,
    \new_Sorter100|1751_ , \new_Sorter100|1752_ , \new_Sorter100|1753_ ,
    \new_Sorter100|1754_ , \new_Sorter100|1755_ , \new_Sorter100|1756_ ,
    \new_Sorter100|1757_ , \new_Sorter100|1758_ , \new_Sorter100|1759_ ,
    \new_Sorter100|1760_ , \new_Sorter100|1761_ , \new_Sorter100|1762_ ,
    \new_Sorter100|1763_ , \new_Sorter100|1764_ , \new_Sorter100|1765_ ,
    \new_Sorter100|1766_ , \new_Sorter100|1767_ , \new_Sorter100|1768_ ,
    \new_Sorter100|1769_ , \new_Sorter100|1770_ , \new_Sorter100|1771_ ,
    \new_Sorter100|1772_ , \new_Sorter100|1773_ , \new_Sorter100|1774_ ,
    \new_Sorter100|1775_ , \new_Sorter100|1776_ , \new_Sorter100|1777_ ,
    \new_Sorter100|1778_ , \new_Sorter100|1779_ , \new_Sorter100|1780_ ,
    \new_Sorter100|1781_ , \new_Sorter100|1782_ , \new_Sorter100|1783_ ,
    \new_Sorter100|1784_ , \new_Sorter100|1785_ , \new_Sorter100|1786_ ,
    \new_Sorter100|1787_ , \new_Sorter100|1788_ , \new_Sorter100|1789_ ,
    \new_Sorter100|1790_ , \new_Sorter100|1791_ , \new_Sorter100|1792_ ,
    \new_Sorter100|1793_ , \new_Sorter100|1794_ , \new_Sorter100|1795_ ,
    \new_Sorter100|1796_ , \new_Sorter100|1797_ , \new_Sorter100|1798_ ,
    \new_Sorter100|1800_ , \new_Sorter100|1801_ , \new_Sorter100|1802_ ,
    \new_Sorter100|1803_ , \new_Sorter100|1804_ , \new_Sorter100|1805_ ,
    \new_Sorter100|1806_ , \new_Sorter100|1807_ , \new_Sorter100|1808_ ,
    \new_Sorter100|1809_ , \new_Sorter100|1810_ , \new_Sorter100|1811_ ,
    \new_Sorter100|1812_ , \new_Sorter100|1813_ , \new_Sorter100|1814_ ,
    \new_Sorter100|1815_ , \new_Sorter100|1816_ , \new_Sorter100|1817_ ,
    \new_Sorter100|1818_ , \new_Sorter100|1819_ , \new_Sorter100|1820_ ,
    \new_Sorter100|1821_ , \new_Sorter100|1822_ , \new_Sorter100|1823_ ,
    \new_Sorter100|1824_ , \new_Sorter100|1825_ , \new_Sorter100|1826_ ,
    \new_Sorter100|1827_ , \new_Sorter100|1828_ , \new_Sorter100|1829_ ,
    \new_Sorter100|1830_ , \new_Sorter100|1831_ , \new_Sorter100|1832_ ,
    \new_Sorter100|1833_ , \new_Sorter100|1834_ , \new_Sorter100|1835_ ,
    \new_Sorter100|1836_ , \new_Sorter100|1837_ , \new_Sorter100|1838_ ,
    \new_Sorter100|1839_ , \new_Sorter100|1840_ , \new_Sorter100|1841_ ,
    \new_Sorter100|1842_ , \new_Sorter100|1843_ , \new_Sorter100|1844_ ,
    \new_Sorter100|1845_ , \new_Sorter100|1846_ , \new_Sorter100|1847_ ,
    \new_Sorter100|1848_ , \new_Sorter100|1849_ , \new_Sorter100|1850_ ,
    \new_Sorter100|1851_ , \new_Sorter100|1852_ , \new_Sorter100|1853_ ,
    \new_Sorter100|1854_ , \new_Sorter100|1855_ , \new_Sorter100|1856_ ,
    \new_Sorter100|1857_ , \new_Sorter100|1858_ , \new_Sorter100|1859_ ,
    \new_Sorter100|1860_ , \new_Sorter100|1861_ , \new_Sorter100|1862_ ,
    \new_Sorter100|1863_ , \new_Sorter100|1864_ , \new_Sorter100|1865_ ,
    \new_Sorter100|1866_ , \new_Sorter100|1867_ , \new_Sorter100|1868_ ,
    \new_Sorter100|1869_ , \new_Sorter100|1870_ , \new_Sorter100|1871_ ,
    \new_Sorter100|1872_ , \new_Sorter100|1873_ , \new_Sorter100|1874_ ,
    \new_Sorter100|1875_ , \new_Sorter100|1876_ , \new_Sorter100|1877_ ,
    \new_Sorter100|1878_ , \new_Sorter100|1879_ , \new_Sorter100|1880_ ,
    \new_Sorter100|1881_ , \new_Sorter100|1882_ , \new_Sorter100|1883_ ,
    \new_Sorter100|1884_ , \new_Sorter100|1885_ , \new_Sorter100|1886_ ,
    \new_Sorter100|1887_ , \new_Sorter100|1888_ , \new_Sorter100|1889_ ,
    \new_Sorter100|1890_ , \new_Sorter100|1891_ , \new_Sorter100|1892_ ,
    \new_Sorter100|1893_ , \new_Sorter100|1894_ , \new_Sorter100|1895_ ,
    \new_Sorter100|1896_ , \new_Sorter100|1897_ , \new_Sorter100|1898_ ,
    \new_Sorter100|1899_ , \new_Sorter100|1900_ , \new_Sorter100|1999_ ,
    \new_Sorter100|1901_ , \new_Sorter100|1902_ , \new_Sorter100|1903_ ,
    \new_Sorter100|1904_ , \new_Sorter100|1905_ , \new_Sorter100|1906_ ,
    \new_Sorter100|1907_ , \new_Sorter100|1908_ , \new_Sorter100|1909_ ,
    \new_Sorter100|1910_ , \new_Sorter100|1911_ , \new_Sorter100|1912_ ,
    \new_Sorter100|1913_ , \new_Sorter100|1914_ , \new_Sorter100|1915_ ,
    \new_Sorter100|1916_ , \new_Sorter100|1917_ , \new_Sorter100|1918_ ,
    \new_Sorter100|1919_ , \new_Sorter100|1920_ , \new_Sorter100|1921_ ,
    \new_Sorter100|1922_ , \new_Sorter100|1923_ , \new_Sorter100|1924_ ,
    \new_Sorter100|1925_ , \new_Sorter100|1926_ , \new_Sorter100|1927_ ,
    \new_Sorter100|1928_ , \new_Sorter100|1929_ , \new_Sorter100|1930_ ,
    \new_Sorter100|1931_ , \new_Sorter100|1932_ , \new_Sorter100|1933_ ,
    \new_Sorter100|1934_ , \new_Sorter100|1935_ , \new_Sorter100|1936_ ,
    \new_Sorter100|1937_ , \new_Sorter100|1938_ , \new_Sorter100|1939_ ,
    \new_Sorter100|1940_ , \new_Sorter100|1941_ , \new_Sorter100|1942_ ,
    \new_Sorter100|1943_ , \new_Sorter100|1944_ , \new_Sorter100|1945_ ,
    \new_Sorter100|1946_ , \new_Sorter100|1947_ , \new_Sorter100|1948_ ,
    \new_Sorter100|1949_ , \new_Sorter100|1950_ , \new_Sorter100|1951_ ,
    \new_Sorter100|1952_ , \new_Sorter100|1953_ , \new_Sorter100|1954_ ,
    \new_Sorter100|1955_ , \new_Sorter100|1956_ , \new_Sorter100|1957_ ,
    \new_Sorter100|1958_ , \new_Sorter100|1959_ , \new_Sorter100|1960_ ,
    \new_Sorter100|1961_ , \new_Sorter100|1962_ , \new_Sorter100|1963_ ,
    \new_Sorter100|1964_ , \new_Sorter100|1965_ , \new_Sorter100|1966_ ,
    \new_Sorter100|1967_ , \new_Sorter100|1968_ , \new_Sorter100|1969_ ,
    \new_Sorter100|1970_ , \new_Sorter100|1971_ , \new_Sorter100|1972_ ,
    \new_Sorter100|1973_ , \new_Sorter100|1974_ , \new_Sorter100|1975_ ,
    \new_Sorter100|1976_ , \new_Sorter100|1977_ , \new_Sorter100|1978_ ,
    \new_Sorter100|1979_ , \new_Sorter100|1980_ , \new_Sorter100|1981_ ,
    \new_Sorter100|1982_ , \new_Sorter100|1983_ , \new_Sorter100|1984_ ,
    \new_Sorter100|1985_ , \new_Sorter100|1986_ , \new_Sorter100|1987_ ,
    \new_Sorter100|1988_ , \new_Sorter100|1989_ , \new_Sorter100|1990_ ,
    \new_Sorter100|1991_ , \new_Sorter100|1992_ , \new_Sorter100|1993_ ,
    \new_Sorter100|1994_ , \new_Sorter100|1995_ , \new_Sorter100|1996_ ,
    \new_Sorter100|1997_ , \new_Sorter100|1998_ , \new_Sorter100|2000_ ,
    \new_Sorter100|2001_ , \new_Sorter100|2002_ , \new_Sorter100|2003_ ,
    \new_Sorter100|2004_ , \new_Sorter100|2005_ , \new_Sorter100|2006_ ,
    \new_Sorter100|2007_ , \new_Sorter100|2008_ , \new_Sorter100|2009_ ,
    \new_Sorter100|2010_ , \new_Sorter100|2011_ , \new_Sorter100|2012_ ,
    \new_Sorter100|2013_ , \new_Sorter100|2014_ , \new_Sorter100|2015_ ,
    \new_Sorter100|2016_ , \new_Sorter100|2017_ , \new_Sorter100|2018_ ,
    \new_Sorter100|2019_ , \new_Sorter100|2020_ , \new_Sorter100|2021_ ,
    \new_Sorter100|2022_ , \new_Sorter100|2023_ , \new_Sorter100|2024_ ,
    \new_Sorter100|2025_ , \new_Sorter100|2026_ , \new_Sorter100|2027_ ,
    \new_Sorter100|2028_ , \new_Sorter100|2029_ , \new_Sorter100|2030_ ,
    \new_Sorter100|2031_ , \new_Sorter100|2032_ , \new_Sorter100|2033_ ,
    \new_Sorter100|2034_ , \new_Sorter100|2035_ , \new_Sorter100|2036_ ,
    \new_Sorter100|2037_ , \new_Sorter100|2038_ , \new_Sorter100|2039_ ,
    \new_Sorter100|2040_ , \new_Sorter100|2041_ , \new_Sorter100|2042_ ,
    \new_Sorter100|2043_ , \new_Sorter100|2044_ , \new_Sorter100|2045_ ,
    \new_Sorter100|2046_ , \new_Sorter100|2047_ , \new_Sorter100|2048_ ,
    \new_Sorter100|2049_ , \new_Sorter100|2050_ , \new_Sorter100|2051_ ,
    \new_Sorter100|2052_ , \new_Sorter100|2053_ , \new_Sorter100|2054_ ,
    \new_Sorter100|2055_ , \new_Sorter100|2056_ , \new_Sorter100|2057_ ,
    \new_Sorter100|2058_ , \new_Sorter100|2059_ , \new_Sorter100|2060_ ,
    \new_Sorter100|2061_ , \new_Sorter100|2062_ , \new_Sorter100|2063_ ,
    \new_Sorter100|2064_ , \new_Sorter100|2065_ , \new_Sorter100|2066_ ,
    \new_Sorter100|2067_ , \new_Sorter100|2068_ , \new_Sorter100|2069_ ,
    \new_Sorter100|2070_ , \new_Sorter100|2071_ , \new_Sorter100|2072_ ,
    \new_Sorter100|2073_ , \new_Sorter100|2074_ , \new_Sorter100|2075_ ,
    \new_Sorter100|2076_ , \new_Sorter100|2077_ , \new_Sorter100|2078_ ,
    \new_Sorter100|2079_ , \new_Sorter100|2080_ , \new_Sorter100|2081_ ,
    \new_Sorter100|2082_ , \new_Sorter100|2083_ , \new_Sorter100|2084_ ,
    \new_Sorter100|2085_ , \new_Sorter100|2086_ , \new_Sorter100|2087_ ,
    \new_Sorter100|2088_ , \new_Sorter100|2089_ , \new_Sorter100|2090_ ,
    \new_Sorter100|2091_ , \new_Sorter100|2092_ , \new_Sorter100|2093_ ,
    \new_Sorter100|2094_ , \new_Sorter100|2095_ , \new_Sorter100|2096_ ,
    \new_Sorter100|2097_ , \new_Sorter100|2098_ , \new_Sorter100|2099_ ,
    \new_Sorter100|2100_ , \new_Sorter100|2199_ , \new_Sorter100|2101_ ,
    \new_Sorter100|2102_ , \new_Sorter100|2103_ , \new_Sorter100|2104_ ,
    \new_Sorter100|2105_ , \new_Sorter100|2106_ , \new_Sorter100|2107_ ,
    \new_Sorter100|2108_ , \new_Sorter100|2109_ , \new_Sorter100|2110_ ,
    \new_Sorter100|2111_ , \new_Sorter100|2112_ , \new_Sorter100|2113_ ,
    \new_Sorter100|2114_ , \new_Sorter100|2115_ , \new_Sorter100|2116_ ,
    \new_Sorter100|2117_ , \new_Sorter100|2118_ , \new_Sorter100|2119_ ,
    \new_Sorter100|2120_ , \new_Sorter100|2121_ , \new_Sorter100|2122_ ,
    \new_Sorter100|2123_ , \new_Sorter100|2124_ , \new_Sorter100|2125_ ,
    \new_Sorter100|2126_ , \new_Sorter100|2127_ , \new_Sorter100|2128_ ,
    \new_Sorter100|2129_ , \new_Sorter100|2130_ , \new_Sorter100|2131_ ,
    \new_Sorter100|2132_ , \new_Sorter100|2133_ , \new_Sorter100|2134_ ,
    \new_Sorter100|2135_ , \new_Sorter100|2136_ , \new_Sorter100|2137_ ,
    \new_Sorter100|2138_ , \new_Sorter100|2139_ , \new_Sorter100|2140_ ,
    \new_Sorter100|2141_ , \new_Sorter100|2142_ , \new_Sorter100|2143_ ,
    \new_Sorter100|2144_ , \new_Sorter100|2145_ , \new_Sorter100|2146_ ,
    \new_Sorter100|2147_ , \new_Sorter100|2148_ , \new_Sorter100|2149_ ,
    \new_Sorter100|2150_ , \new_Sorter100|2151_ , \new_Sorter100|2152_ ,
    \new_Sorter100|2153_ , \new_Sorter100|2154_ , \new_Sorter100|2155_ ,
    \new_Sorter100|2156_ , \new_Sorter100|2157_ , \new_Sorter100|2158_ ,
    \new_Sorter100|2159_ , \new_Sorter100|2160_ , \new_Sorter100|2161_ ,
    \new_Sorter100|2162_ , \new_Sorter100|2163_ , \new_Sorter100|2164_ ,
    \new_Sorter100|2165_ , \new_Sorter100|2166_ , \new_Sorter100|2167_ ,
    \new_Sorter100|2168_ , \new_Sorter100|2169_ , \new_Sorter100|2170_ ,
    \new_Sorter100|2171_ , \new_Sorter100|2172_ , \new_Sorter100|2173_ ,
    \new_Sorter100|2174_ , \new_Sorter100|2175_ , \new_Sorter100|2176_ ,
    \new_Sorter100|2177_ , \new_Sorter100|2178_ , \new_Sorter100|2179_ ,
    \new_Sorter100|2180_ , \new_Sorter100|2181_ , \new_Sorter100|2182_ ,
    \new_Sorter100|2183_ , \new_Sorter100|2184_ , \new_Sorter100|2185_ ,
    \new_Sorter100|2186_ , \new_Sorter100|2187_ , \new_Sorter100|2188_ ,
    \new_Sorter100|2189_ , \new_Sorter100|2190_ , \new_Sorter100|2191_ ,
    \new_Sorter100|2192_ , \new_Sorter100|2193_ , \new_Sorter100|2194_ ,
    \new_Sorter100|2195_ , \new_Sorter100|2196_ , \new_Sorter100|2197_ ,
    \new_Sorter100|2198_ , \new_Sorter100|2200_ , \new_Sorter100|2201_ ,
    \new_Sorter100|2202_ , \new_Sorter100|2203_ , \new_Sorter100|2204_ ,
    \new_Sorter100|2205_ , \new_Sorter100|2206_ , \new_Sorter100|2207_ ,
    \new_Sorter100|2208_ , \new_Sorter100|2209_ , \new_Sorter100|2210_ ,
    \new_Sorter100|2211_ , \new_Sorter100|2212_ , \new_Sorter100|2213_ ,
    \new_Sorter100|2214_ , \new_Sorter100|2215_ , \new_Sorter100|2216_ ,
    \new_Sorter100|2217_ , \new_Sorter100|2218_ , \new_Sorter100|2219_ ,
    \new_Sorter100|2220_ , \new_Sorter100|2221_ , \new_Sorter100|2222_ ,
    \new_Sorter100|2223_ , \new_Sorter100|2224_ , \new_Sorter100|2225_ ,
    \new_Sorter100|2226_ , \new_Sorter100|2227_ , \new_Sorter100|2228_ ,
    \new_Sorter100|2229_ , \new_Sorter100|2230_ , \new_Sorter100|2231_ ,
    \new_Sorter100|2232_ , \new_Sorter100|2233_ , \new_Sorter100|2234_ ,
    \new_Sorter100|2235_ , \new_Sorter100|2236_ , \new_Sorter100|2237_ ,
    \new_Sorter100|2238_ , \new_Sorter100|2239_ , \new_Sorter100|2240_ ,
    \new_Sorter100|2241_ , \new_Sorter100|2242_ , \new_Sorter100|2243_ ,
    \new_Sorter100|2244_ , \new_Sorter100|2245_ , \new_Sorter100|2246_ ,
    \new_Sorter100|2247_ , \new_Sorter100|2248_ , \new_Sorter100|2249_ ,
    \new_Sorter100|2250_ , \new_Sorter100|2251_ , \new_Sorter100|2252_ ,
    \new_Sorter100|2253_ , \new_Sorter100|2254_ , \new_Sorter100|2255_ ,
    \new_Sorter100|2256_ , \new_Sorter100|2257_ , \new_Sorter100|2258_ ,
    \new_Sorter100|2259_ , \new_Sorter100|2260_ , \new_Sorter100|2261_ ,
    \new_Sorter100|2262_ , \new_Sorter100|2263_ , \new_Sorter100|2264_ ,
    \new_Sorter100|2265_ , \new_Sorter100|2266_ , \new_Sorter100|2267_ ,
    \new_Sorter100|2268_ , \new_Sorter100|2269_ , \new_Sorter100|2270_ ,
    \new_Sorter100|2271_ , \new_Sorter100|2272_ , \new_Sorter100|2273_ ,
    \new_Sorter100|2274_ , \new_Sorter100|2275_ , \new_Sorter100|2276_ ,
    \new_Sorter100|2277_ , \new_Sorter100|2278_ , \new_Sorter100|2279_ ,
    \new_Sorter100|2280_ , \new_Sorter100|2281_ , \new_Sorter100|2282_ ,
    \new_Sorter100|2283_ , \new_Sorter100|2284_ , \new_Sorter100|2285_ ,
    \new_Sorter100|2286_ , \new_Sorter100|2287_ , \new_Sorter100|2288_ ,
    \new_Sorter100|2289_ , \new_Sorter100|2290_ , \new_Sorter100|2291_ ,
    \new_Sorter100|2292_ , \new_Sorter100|2293_ , \new_Sorter100|2294_ ,
    \new_Sorter100|2295_ , \new_Sorter100|2296_ , \new_Sorter100|2297_ ,
    \new_Sorter100|2298_ , \new_Sorter100|2299_ , \new_Sorter100|2300_ ,
    \new_Sorter100|2399_ , \new_Sorter100|2301_ , \new_Sorter100|2302_ ,
    \new_Sorter100|2303_ , \new_Sorter100|2304_ , \new_Sorter100|2305_ ,
    \new_Sorter100|2306_ , \new_Sorter100|2307_ , \new_Sorter100|2308_ ,
    \new_Sorter100|2309_ , \new_Sorter100|2310_ , \new_Sorter100|2311_ ,
    \new_Sorter100|2312_ , \new_Sorter100|2313_ , \new_Sorter100|2314_ ,
    \new_Sorter100|2315_ , \new_Sorter100|2316_ , \new_Sorter100|2317_ ,
    \new_Sorter100|2318_ , \new_Sorter100|2319_ , \new_Sorter100|2320_ ,
    \new_Sorter100|2321_ , \new_Sorter100|2322_ , \new_Sorter100|2323_ ,
    \new_Sorter100|2324_ , \new_Sorter100|2325_ , \new_Sorter100|2326_ ,
    \new_Sorter100|2327_ , \new_Sorter100|2328_ , \new_Sorter100|2329_ ,
    \new_Sorter100|2330_ , \new_Sorter100|2331_ , \new_Sorter100|2332_ ,
    \new_Sorter100|2333_ , \new_Sorter100|2334_ , \new_Sorter100|2335_ ,
    \new_Sorter100|2336_ , \new_Sorter100|2337_ , \new_Sorter100|2338_ ,
    \new_Sorter100|2339_ , \new_Sorter100|2340_ , \new_Sorter100|2341_ ,
    \new_Sorter100|2342_ , \new_Sorter100|2343_ , \new_Sorter100|2344_ ,
    \new_Sorter100|2345_ , \new_Sorter100|2346_ , \new_Sorter100|2347_ ,
    \new_Sorter100|2348_ , \new_Sorter100|2349_ , \new_Sorter100|2350_ ,
    \new_Sorter100|2351_ , \new_Sorter100|2352_ , \new_Sorter100|2353_ ,
    \new_Sorter100|2354_ , \new_Sorter100|2355_ , \new_Sorter100|2356_ ,
    \new_Sorter100|2357_ , \new_Sorter100|2358_ , \new_Sorter100|2359_ ,
    \new_Sorter100|2360_ , \new_Sorter100|2361_ , \new_Sorter100|2362_ ,
    \new_Sorter100|2363_ , \new_Sorter100|2364_ , \new_Sorter100|2365_ ,
    \new_Sorter100|2366_ , \new_Sorter100|2367_ , \new_Sorter100|2368_ ,
    \new_Sorter100|2369_ , \new_Sorter100|2370_ , \new_Sorter100|2371_ ,
    \new_Sorter100|2372_ , \new_Sorter100|2373_ , \new_Sorter100|2374_ ,
    \new_Sorter100|2375_ , \new_Sorter100|2376_ , \new_Sorter100|2377_ ,
    \new_Sorter100|2378_ , \new_Sorter100|2379_ , \new_Sorter100|2380_ ,
    \new_Sorter100|2381_ , \new_Sorter100|2382_ , \new_Sorter100|2383_ ,
    \new_Sorter100|2384_ , \new_Sorter100|2385_ , \new_Sorter100|2386_ ,
    \new_Sorter100|2387_ , \new_Sorter100|2388_ , \new_Sorter100|2389_ ,
    \new_Sorter100|2390_ , \new_Sorter100|2391_ , \new_Sorter100|2392_ ,
    \new_Sorter100|2393_ , \new_Sorter100|2394_ , \new_Sorter100|2395_ ,
    \new_Sorter100|2396_ , \new_Sorter100|2397_ , \new_Sorter100|2398_ ,
    \new_Sorter100|2400_ , \new_Sorter100|2401_ , \new_Sorter100|2402_ ,
    \new_Sorter100|2403_ , \new_Sorter100|2404_ , \new_Sorter100|2405_ ,
    \new_Sorter100|2406_ , \new_Sorter100|2407_ , \new_Sorter100|2408_ ,
    \new_Sorter100|2409_ , \new_Sorter100|2410_ , \new_Sorter100|2411_ ,
    \new_Sorter100|2412_ , \new_Sorter100|2413_ , \new_Sorter100|2414_ ,
    \new_Sorter100|2415_ , \new_Sorter100|2416_ , \new_Sorter100|2417_ ,
    \new_Sorter100|2418_ , \new_Sorter100|2419_ , \new_Sorter100|2420_ ,
    \new_Sorter100|2421_ , \new_Sorter100|2422_ , \new_Sorter100|2423_ ,
    \new_Sorter100|2424_ , \new_Sorter100|2425_ , \new_Sorter100|2426_ ,
    \new_Sorter100|2427_ , \new_Sorter100|2428_ , \new_Sorter100|2429_ ,
    \new_Sorter100|2430_ , \new_Sorter100|2431_ , \new_Sorter100|2432_ ,
    \new_Sorter100|2433_ , \new_Sorter100|2434_ , \new_Sorter100|2435_ ,
    \new_Sorter100|2436_ , \new_Sorter100|2437_ , \new_Sorter100|2438_ ,
    \new_Sorter100|2439_ , \new_Sorter100|2440_ , \new_Sorter100|2441_ ,
    \new_Sorter100|2442_ , \new_Sorter100|2443_ , \new_Sorter100|2444_ ,
    \new_Sorter100|2445_ , \new_Sorter100|2446_ , \new_Sorter100|2447_ ,
    \new_Sorter100|2448_ , \new_Sorter100|2449_ , \new_Sorter100|2450_ ,
    \new_Sorter100|2451_ , \new_Sorter100|2452_ , \new_Sorter100|2453_ ,
    \new_Sorter100|2454_ , \new_Sorter100|2455_ , \new_Sorter100|2456_ ,
    \new_Sorter100|2457_ , \new_Sorter100|2458_ , \new_Sorter100|2459_ ,
    \new_Sorter100|2460_ , \new_Sorter100|2461_ , \new_Sorter100|2462_ ,
    \new_Sorter100|2463_ , \new_Sorter100|2464_ , \new_Sorter100|2465_ ,
    \new_Sorter100|2466_ , \new_Sorter100|2467_ , \new_Sorter100|2468_ ,
    \new_Sorter100|2469_ , \new_Sorter100|2470_ , \new_Sorter100|2471_ ,
    \new_Sorter100|2472_ , \new_Sorter100|2473_ , \new_Sorter100|2474_ ,
    \new_Sorter100|2475_ , \new_Sorter100|2476_ , \new_Sorter100|2477_ ,
    \new_Sorter100|2478_ , \new_Sorter100|2479_ , \new_Sorter100|2480_ ,
    \new_Sorter100|2481_ , \new_Sorter100|2482_ , \new_Sorter100|2483_ ,
    \new_Sorter100|2484_ , \new_Sorter100|2485_ , \new_Sorter100|2486_ ,
    \new_Sorter100|2487_ , \new_Sorter100|2488_ , \new_Sorter100|2489_ ,
    \new_Sorter100|2490_ , \new_Sorter100|2491_ , \new_Sorter100|2492_ ,
    \new_Sorter100|2493_ , \new_Sorter100|2494_ , \new_Sorter100|2495_ ,
    \new_Sorter100|2496_ , \new_Sorter100|2497_ , \new_Sorter100|2498_ ,
    \new_Sorter100|2499_ , \new_Sorter100|2500_ , \new_Sorter100|2599_ ,
    \new_Sorter100|2501_ , \new_Sorter100|2502_ , \new_Sorter100|2503_ ,
    \new_Sorter100|2504_ , \new_Sorter100|2505_ , \new_Sorter100|2506_ ,
    \new_Sorter100|2507_ , \new_Sorter100|2508_ , \new_Sorter100|2509_ ,
    \new_Sorter100|2510_ , \new_Sorter100|2511_ , \new_Sorter100|2512_ ,
    \new_Sorter100|2513_ , \new_Sorter100|2514_ , \new_Sorter100|2515_ ,
    \new_Sorter100|2516_ , \new_Sorter100|2517_ , \new_Sorter100|2518_ ,
    \new_Sorter100|2519_ , \new_Sorter100|2520_ , \new_Sorter100|2521_ ,
    \new_Sorter100|2522_ , \new_Sorter100|2523_ , \new_Sorter100|2524_ ,
    \new_Sorter100|2525_ , \new_Sorter100|2526_ , \new_Sorter100|2527_ ,
    \new_Sorter100|2528_ , \new_Sorter100|2529_ , \new_Sorter100|2530_ ,
    \new_Sorter100|2531_ , \new_Sorter100|2532_ , \new_Sorter100|2533_ ,
    \new_Sorter100|2534_ , \new_Sorter100|2535_ , \new_Sorter100|2536_ ,
    \new_Sorter100|2537_ , \new_Sorter100|2538_ , \new_Sorter100|2539_ ,
    \new_Sorter100|2540_ , \new_Sorter100|2541_ , \new_Sorter100|2542_ ,
    \new_Sorter100|2543_ , \new_Sorter100|2544_ , \new_Sorter100|2545_ ,
    \new_Sorter100|2546_ , \new_Sorter100|2547_ , \new_Sorter100|2548_ ,
    \new_Sorter100|2549_ , \new_Sorter100|2550_ , \new_Sorter100|2551_ ,
    \new_Sorter100|2552_ , \new_Sorter100|2553_ , \new_Sorter100|2554_ ,
    \new_Sorter100|2555_ , \new_Sorter100|2556_ , \new_Sorter100|2557_ ,
    \new_Sorter100|2558_ , \new_Sorter100|2559_ , \new_Sorter100|2560_ ,
    \new_Sorter100|2561_ , \new_Sorter100|2562_ , \new_Sorter100|2563_ ,
    \new_Sorter100|2564_ , \new_Sorter100|2565_ , \new_Sorter100|2566_ ,
    \new_Sorter100|2567_ , \new_Sorter100|2568_ , \new_Sorter100|2569_ ,
    \new_Sorter100|2570_ , \new_Sorter100|2571_ , \new_Sorter100|2572_ ,
    \new_Sorter100|2573_ , \new_Sorter100|2574_ , \new_Sorter100|2575_ ,
    \new_Sorter100|2576_ , \new_Sorter100|2577_ , \new_Sorter100|2578_ ,
    \new_Sorter100|2579_ , \new_Sorter100|2580_ , \new_Sorter100|2581_ ,
    \new_Sorter100|2582_ , \new_Sorter100|2583_ , \new_Sorter100|2584_ ,
    \new_Sorter100|2585_ , \new_Sorter100|2586_ , \new_Sorter100|2587_ ,
    \new_Sorter100|2588_ , \new_Sorter100|2589_ , \new_Sorter100|2590_ ,
    \new_Sorter100|2591_ , \new_Sorter100|2592_ , \new_Sorter100|2593_ ,
    \new_Sorter100|2594_ , \new_Sorter100|2595_ , \new_Sorter100|2596_ ,
    \new_Sorter100|2597_ , \new_Sorter100|2598_ , \new_Sorter100|2600_ ,
    \new_Sorter100|2601_ , \new_Sorter100|2602_ , \new_Sorter100|2603_ ,
    \new_Sorter100|2604_ , \new_Sorter100|2605_ , \new_Sorter100|2606_ ,
    \new_Sorter100|2607_ , \new_Sorter100|2608_ , \new_Sorter100|2609_ ,
    \new_Sorter100|2610_ , \new_Sorter100|2611_ , \new_Sorter100|2612_ ,
    \new_Sorter100|2613_ , \new_Sorter100|2614_ , \new_Sorter100|2615_ ,
    \new_Sorter100|2616_ , \new_Sorter100|2617_ , \new_Sorter100|2618_ ,
    \new_Sorter100|2619_ , \new_Sorter100|2620_ , \new_Sorter100|2621_ ,
    \new_Sorter100|2622_ , \new_Sorter100|2623_ , \new_Sorter100|2624_ ,
    \new_Sorter100|2625_ , \new_Sorter100|2626_ , \new_Sorter100|2627_ ,
    \new_Sorter100|2628_ , \new_Sorter100|2629_ , \new_Sorter100|2630_ ,
    \new_Sorter100|2631_ , \new_Sorter100|2632_ , \new_Sorter100|2633_ ,
    \new_Sorter100|2634_ , \new_Sorter100|2635_ , \new_Sorter100|2636_ ,
    \new_Sorter100|2637_ , \new_Sorter100|2638_ , \new_Sorter100|2639_ ,
    \new_Sorter100|2640_ , \new_Sorter100|2641_ , \new_Sorter100|2642_ ,
    \new_Sorter100|2643_ , \new_Sorter100|2644_ , \new_Sorter100|2645_ ,
    \new_Sorter100|2646_ , \new_Sorter100|2647_ , \new_Sorter100|2648_ ,
    \new_Sorter100|2649_ , \new_Sorter100|2650_ , \new_Sorter100|2651_ ,
    \new_Sorter100|2652_ , \new_Sorter100|2653_ , \new_Sorter100|2654_ ,
    \new_Sorter100|2655_ , \new_Sorter100|2656_ , \new_Sorter100|2657_ ,
    \new_Sorter100|2658_ , \new_Sorter100|2659_ , \new_Sorter100|2660_ ,
    \new_Sorter100|2661_ , \new_Sorter100|2662_ , \new_Sorter100|2663_ ,
    \new_Sorter100|2664_ , \new_Sorter100|2665_ , \new_Sorter100|2666_ ,
    \new_Sorter100|2667_ , \new_Sorter100|2668_ , \new_Sorter100|2669_ ,
    \new_Sorter100|2670_ , \new_Sorter100|2671_ , \new_Sorter100|2672_ ,
    \new_Sorter100|2673_ , \new_Sorter100|2674_ , \new_Sorter100|2675_ ,
    \new_Sorter100|2676_ , \new_Sorter100|2677_ , \new_Sorter100|2678_ ,
    \new_Sorter100|2679_ , \new_Sorter100|2680_ , \new_Sorter100|2681_ ,
    \new_Sorter100|2682_ , \new_Sorter100|2683_ , \new_Sorter100|2684_ ,
    \new_Sorter100|2685_ , \new_Sorter100|2686_ , \new_Sorter100|2687_ ,
    \new_Sorter100|2688_ , \new_Sorter100|2689_ , \new_Sorter100|2690_ ,
    \new_Sorter100|2691_ , \new_Sorter100|2692_ , \new_Sorter100|2693_ ,
    \new_Sorter100|2694_ , \new_Sorter100|2695_ , \new_Sorter100|2696_ ,
    \new_Sorter100|2697_ , \new_Sorter100|2698_ , \new_Sorter100|2699_ ,
    \new_Sorter100|2700_ , \new_Sorter100|2799_ , \new_Sorter100|2701_ ,
    \new_Sorter100|2702_ , \new_Sorter100|2703_ , \new_Sorter100|2704_ ,
    \new_Sorter100|2705_ , \new_Sorter100|2706_ , \new_Sorter100|2707_ ,
    \new_Sorter100|2708_ , \new_Sorter100|2709_ , \new_Sorter100|2710_ ,
    \new_Sorter100|2711_ , \new_Sorter100|2712_ , \new_Sorter100|2713_ ,
    \new_Sorter100|2714_ , \new_Sorter100|2715_ , \new_Sorter100|2716_ ,
    \new_Sorter100|2717_ , \new_Sorter100|2718_ , \new_Sorter100|2719_ ,
    \new_Sorter100|2720_ , \new_Sorter100|2721_ , \new_Sorter100|2722_ ,
    \new_Sorter100|2723_ , \new_Sorter100|2724_ , \new_Sorter100|2725_ ,
    \new_Sorter100|2726_ , \new_Sorter100|2727_ , \new_Sorter100|2728_ ,
    \new_Sorter100|2729_ , \new_Sorter100|2730_ , \new_Sorter100|2731_ ,
    \new_Sorter100|2732_ , \new_Sorter100|2733_ , \new_Sorter100|2734_ ,
    \new_Sorter100|2735_ , \new_Sorter100|2736_ , \new_Sorter100|2737_ ,
    \new_Sorter100|2738_ , \new_Sorter100|2739_ , \new_Sorter100|2740_ ,
    \new_Sorter100|2741_ , \new_Sorter100|2742_ , \new_Sorter100|2743_ ,
    \new_Sorter100|2744_ , \new_Sorter100|2745_ , \new_Sorter100|2746_ ,
    \new_Sorter100|2747_ , \new_Sorter100|2748_ , \new_Sorter100|2749_ ,
    \new_Sorter100|2750_ , \new_Sorter100|2751_ , \new_Sorter100|2752_ ,
    \new_Sorter100|2753_ , \new_Sorter100|2754_ , \new_Sorter100|2755_ ,
    \new_Sorter100|2756_ , \new_Sorter100|2757_ , \new_Sorter100|2758_ ,
    \new_Sorter100|2759_ , \new_Sorter100|2760_ , \new_Sorter100|2761_ ,
    \new_Sorter100|2762_ , \new_Sorter100|2763_ , \new_Sorter100|2764_ ,
    \new_Sorter100|2765_ , \new_Sorter100|2766_ , \new_Sorter100|2767_ ,
    \new_Sorter100|2768_ , \new_Sorter100|2769_ , \new_Sorter100|2770_ ,
    \new_Sorter100|2771_ , \new_Sorter100|2772_ , \new_Sorter100|2773_ ,
    \new_Sorter100|2774_ , \new_Sorter100|2775_ , \new_Sorter100|2776_ ,
    \new_Sorter100|2777_ , \new_Sorter100|2778_ , \new_Sorter100|2779_ ,
    \new_Sorter100|2780_ , \new_Sorter100|2781_ , \new_Sorter100|2782_ ,
    \new_Sorter100|2783_ , \new_Sorter100|2784_ , \new_Sorter100|2785_ ,
    \new_Sorter100|2786_ , \new_Sorter100|2787_ , \new_Sorter100|2788_ ,
    \new_Sorter100|2789_ , \new_Sorter100|2790_ , \new_Sorter100|2791_ ,
    \new_Sorter100|2792_ , \new_Sorter100|2793_ , \new_Sorter100|2794_ ,
    \new_Sorter100|2795_ , \new_Sorter100|2796_ , \new_Sorter100|2797_ ,
    \new_Sorter100|2798_ , \new_Sorter100|2800_ , \new_Sorter100|2801_ ,
    \new_Sorter100|2802_ , \new_Sorter100|2803_ , \new_Sorter100|2804_ ,
    \new_Sorter100|2805_ , \new_Sorter100|2806_ , \new_Sorter100|2807_ ,
    \new_Sorter100|2808_ , \new_Sorter100|2809_ , \new_Sorter100|2810_ ,
    \new_Sorter100|2811_ , \new_Sorter100|2812_ , \new_Sorter100|2813_ ,
    \new_Sorter100|2814_ , \new_Sorter100|2815_ , \new_Sorter100|2816_ ,
    \new_Sorter100|2817_ , \new_Sorter100|2818_ , \new_Sorter100|2819_ ,
    \new_Sorter100|2820_ , \new_Sorter100|2821_ , \new_Sorter100|2822_ ,
    \new_Sorter100|2823_ , \new_Sorter100|2824_ , \new_Sorter100|2825_ ,
    \new_Sorter100|2826_ , \new_Sorter100|2827_ , \new_Sorter100|2828_ ,
    \new_Sorter100|2829_ , \new_Sorter100|2830_ , \new_Sorter100|2831_ ,
    \new_Sorter100|2832_ , \new_Sorter100|2833_ , \new_Sorter100|2834_ ,
    \new_Sorter100|2835_ , \new_Sorter100|2836_ , \new_Sorter100|2837_ ,
    \new_Sorter100|2838_ , \new_Sorter100|2839_ , \new_Sorter100|2840_ ,
    \new_Sorter100|2841_ , \new_Sorter100|2842_ , \new_Sorter100|2843_ ,
    \new_Sorter100|2844_ , \new_Sorter100|2845_ , \new_Sorter100|2846_ ,
    \new_Sorter100|2847_ , \new_Sorter100|2848_ , \new_Sorter100|2849_ ,
    \new_Sorter100|2850_ , \new_Sorter100|2851_ , \new_Sorter100|2852_ ,
    \new_Sorter100|2853_ , \new_Sorter100|2854_ , \new_Sorter100|2855_ ,
    \new_Sorter100|2856_ , \new_Sorter100|2857_ , \new_Sorter100|2858_ ,
    \new_Sorter100|2859_ , \new_Sorter100|2860_ , \new_Sorter100|2861_ ,
    \new_Sorter100|2862_ , \new_Sorter100|2863_ , \new_Sorter100|2864_ ,
    \new_Sorter100|2865_ , \new_Sorter100|2866_ , \new_Sorter100|2867_ ,
    \new_Sorter100|2868_ , \new_Sorter100|2869_ , \new_Sorter100|2870_ ,
    \new_Sorter100|2871_ , \new_Sorter100|2872_ , \new_Sorter100|2873_ ,
    \new_Sorter100|2874_ , \new_Sorter100|2875_ , \new_Sorter100|2876_ ,
    \new_Sorter100|2877_ , \new_Sorter100|2878_ , \new_Sorter100|2879_ ,
    \new_Sorter100|2880_ , \new_Sorter100|2881_ , \new_Sorter100|2882_ ,
    \new_Sorter100|2883_ , \new_Sorter100|2884_ , \new_Sorter100|2885_ ,
    \new_Sorter100|2886_ , \new_Sorter100|2887_ , \new_Sorter100|2888_ ,
    \new_Sorter100|2889_ , \new_Sorter100|2890_ , \new_Sorter100|2891_ ,
    \new_Sorter100|2892_ , \new_Sorter100|2893_ , \new_Sorter100|2894_ ,
    \new_Sorter100|2895_ , \new_Sorter100|2896_ , \new_Sorter100|2897_ ,
    \new_Sorter100|2898_ , \new_Sorter100|2899_ , \new_Sorter100|2900_ ,
    \new_Sorter100|2999_ , \new_Sorter100|2901_ , \new_Sorter100|2902_ ,
    \new_Sorter100|2903_ , \new_Sorter100|2904_ , \new_Sorter100|2905_ ,
    \new_Sorter100|2906_ , \new_Sorter100|2907_ , \new_Sorter100|2908_ ,
    \new_Sorter100|2909_ , \new_Sorter100|2910_ , \new_Sorter100|2911_ ,
    \new_Sorter100|2912_ , \new_Sorter100|2913_ , \new_Sorter100|2914_ ,
    \new_Sorter100|2915_ , \new_Sorter100|2916_ , \new_Sorter100|2917_ ,
    \new_Sorter100|2918_ , \new_Sorter100|2919_ , \new_Sorter100|2920_ ,
    \new_Sorter100|2921_ , \new_Sorter100|2922_ , \new_Sorter100|2923_ ,
    \new_Sorter100|2924_ , \new_Sorter100|2925_ , \new_Sorter100|2926_ ,
    \new_Sorter100|2927_ , \new_Sorter100|2928_ , \new_Sorter100|2929_ ,
    \new_Sorter100|2930_ , \new_Sorter100|2931_ , \new_Sorter100|2932_ ,
    \new_Sorter100|2933_ , \new_Sorter100|2934_ , \new_Sorter100|2935_ ,
    \new_Sorter100|2936_ , \new_Sorter100|2937_ , \new_Sorter100|2938_ ,
    \new_Sorter100|2939_ , \new_Sorter100|2940_ , \new_Sorter100|2941_ ,
    \new_Sorter100|2942_ , \new_Sorter100|2943_ , \new_Sorter100|2944_ ,
    \new_Sorter100|2945_ , \new_Sorter100|2946_ , \new_Sorter100|2947_ ,
    \new_Sorter100|2948_ , \new_Sorter100|2949_ , \new_Sorter100|2950_ ,
    \new_Sorter100|2951_ , \new_Sorter100|2952_ , \new_Sorter100|2953_ ,
    \new_Sorter100|2954_ , \new_Sorter100|2955_ , \new_Sorter100|2956_ ,
    \new_Sorter100|2957_ , \new_Sorter100|2958_ , \new_Sorter100|2959_ ,
    \new_Sorter100|2960_ , \new_Sorter100|2961_ , \new_Sorter100|2962_ ,
    \new_Sorter100|2963_ , \new_Sorter100|2964_ , \new_Sorter100|2965_ ,
    \new_Sorter100|2966_ , \new_Sorter100|2967_ , \new_Sorter100|2968_ ,
    \new_Sorter100|2969_ , \new_Sorter100|2970_ , \new_Sorter100|2971_ ,
    \new_Sorter100|2972_ , \new_Sorter100|2973_ , \new_Sorter100|2974_ ,
    \new_Sorter100|2975_ , \new_Sorter100|2976_ , \new_Sorter100|2977_ ,
    \new_Sorter100|2978_ , \new_Sorter100|2979_ , \new_Sorter100|2980_ ,
    \new_Sorter100|2981_ , \new_Sorter100|2982_ , \new_Sorter100|2983_ ,
    \new_Sorter100|2984_ , \new_Sorter100|2985_ , \new_Sorter100|2986_ ,
    \new_Sorter100|2987_ , \new_Sorter100|2988_ , \new_Sorter100|2989_ ,
    \new_Sorter100|2990_ , \new_Sorter100|2991_ , \new_Sorter100|2992_ ,
    \new_Sorter100|2993_ , \new_Sorter100|2994_ , \new_Sorter100|2995_ ,
    \new_Sorter100|2996_ , \new_Sorter100|2997_ , \new_Sorter100|2998_ ,
    \new_Sorter100|3000_ , \new_Sorter100|3001_ , \new_Sorter100|3002_ ,
    \new_Sorter100|3003_ , \new_Sorter100|3004_ , \new_Sorter100|3005_ ,
    \new_Sorter100|3006_ , \new_Sorter100|3007_ , \new_Sorter100|3008_ ,
    \new_Sorter100|3009_ , \new_Sorter100|3010_ , \new_Sorter100|3011_ ,
    \new_Sorter100|3012_ , \new_Sorter100|3013_ , \new_Sorter100|3014_ ,
    \new_Sorter100|3015_ , \new_Sorter100|3016_ , \new_Sorter100|3017_ ,
    \new_Sorter100|3018_ , \new_Sorter100|3019_ , \new_Sorter100|3020_ ,
    \new_Sorter100|3021_ , \new_Sorter100|3022_ , \new_Sorter100|3023_ ,
    \new_Sorter100|3024_ , \new_Sorter100|3025_ , \new_Sorter100|3026_ ,
    \new_Sorter100|3027_ , \new_Sorter100|3028_ , \new_Sorter100|3029_ ,
    \new_Sorter100|3030_ , \new_Sorter100|3031_ , \new_Sorter100|3032_ ,
    \new_Sorter100|3033_ , \new_Sorter100|3034_ , \new_Sorter100|3035_ ,
    \new_Sorter100|3036_ , \new_Sorter100|3037_ , \new_Sorter100|3038_ ,
    \new_Sorter100|3039_ , \new_Sorter100|3040_ , \new_Sorter100|3041_ ,
    \new_Sorter100|3042_ , \new_Sorter100|3043_ , \new_Sorter100|3044_ ,
    \new_Sorter100|3045_ , \new_Sorter100|3046_ , \new_Sorter100|3047_ ,
    \new_Sorter100|3048_ , \new_Sorter100|3049_ , \new_Sorter100|3050_ ,
    \new_Sorter100|3051_ , \new_Sorter100|3052_ , \new_Sorter100|3053_ ,
    \new_Sorter100|3054_ , \new_Sorter100|3055_ , \new_Sorter100|3056_ ,
    \new_Sorter100|3057_ , \new_Sorter100|3058_ , \new_Sorter100|3059_ ,
    \new_Sorter100|3060_ , \new_Sorter100|3061_ , \new_Sorter100|3062_ ,
    \new_Sorter100|3063_ , \new_Sorter100|3064_ , \new_Sorter100|3065_ ,
    \new_Sorter100|3066_ , \new_Sorter100|3067_ , \new_Sorter100|3068_ ,
    \new_Sorter100|3069_ , \new_Sorter100|3070_ , \new_Sorter100|3071_ ,
    \new_Sorter100|3072_ , \new_Sorter100|3073_ , \new_Sorter100|3074_ ,
    \new_Sorter100|3075_ , \new_Sorter100|3076_ , \new_Sorter100|3077_ ,
    \new_Sorter100|3078_ , \new_Sorter100|3079_ , \new_Sorter100|3080_ ,
    \new_Sorter100|3081_ , \new_Sorter100|3082_ , \new_Sorter100|3083_ ,
    \new_Sorter100|3084_ , \new_Sorter100|3085_ , \new_Sorter100|3086_ ,
    \new_Sorter100|3087_ , \new_Sorter100|3088_ , \new_Sorter100|3089_ ,
    \new_Sorter100|3090_ , \new_Sorter100|3091_ , \new_Sorter100|3092_ ,
    \new_Sorter100|3093_ , \new_Sorter100|3094_ , \new_Sorter100|3095_ ,
    \new_Sorter100|3096_ , \new_Sorter100|3097_ , \new_Sorter100|3098_ ,
    \new_Sorter100|3099_ , \new_Sorter100|3100_ , \new_Sorter100|3199_ ,
    \new_Sorter100|3101_ , \new_Sorter100|3102_ , \new_Sorter100|3103_ ,
    \new_Sorter100|3104_ , \new_Sorter100|3105_ , \new_Sorter100|3106_ ,
    \new_Sorter100|3107_ , \new_Sorter100|3108_ , \new_Sorter100|3109_ ,
    \new_Sorter100|3110_ , \new_Sorter100|3111_ , \new_Sorter100|3112_ ,
    \new_Sorter100|3113_ , \new_Sorter100|3114_ , \new_Sorter100|3115_ ,
    \new_Sorter100|3116_ , \new_Sorter100|3117_ , \new_Sorter100|3118_ ,
    \new_Sorter100|3119_ , \new_Sorter100|3120_ , \new_Sorter100|3121_ ,
    \new_Sorter100|3122_ , \new_Sorter100|3123_ , \new_Sorter100|3124_ ,
    \new_Sorter100|3125_ , \new_Sorter100|3126_ , \new_Sorter100|3127_ ,
    \new_Sorter100|3128_ , \new_Sorter100|3129_ , \new_Sorter100|3130_ ,
    \new_Sorter100|3131_ , \new_Sorter100|3132_ , \new_Sorter100|3133_ ,
    \new_Sorter100|3134_ , \new_Sorter100|3135_ , \new_Sorter100|3136_ ,
    \new_Sorter100|3137_ , \new_Sorter100|3138_ , \new_Sorter100|3139_ ,
    \new_Sorter100|3140_ , \new_Sorter100|3141_ , \new_Sorter100|3142_ ,
    \new_Sorter100|3143_ , \new_Sorter100|3144_ , \new_Sorter100|3145_ ,
    \new_Sorter100|3146_ , \new_Sorter100|3147_ , \new_Sorter100|3148_ ,
    \new_Sorter100|3149_ , \new_Sorter100|3150_ , \new_Sorter100|3151_ ,
    \new_Sorter100|3152_ , \new_Sorter100|3153_ , \new_Sorter100|3154_ ,
    \new_Sorter100|3155_ , \new_Sorter100|3156_ , \new_Sorter100|3157_ ,
    \new_Sorter100|3158_ , \new_Sorter100|3159_ , \new_Sorter100|3160_ ,
    \new_Sorter100|3161_ , \new_Sorter100|3162_ , \new_Sorter100|3163_ ,
    \new_Sorter100|3164_ , \new_Sorter100|3165_ , \new_Sorter100|3166_ ,
    \new_Sorter100|3167_ , \new_Sorter100|3168_ , \new_Sorter100|3169_ ,
    \new_Sorter100|3170_ , \new_Sorter100|3171_ , \new_Sorter100|3172_ ,
    \new_Sorter100|3173_ , \new_Sorter100|3174_ , \new_Sorter100|3175_ ,
    \new_Sorter100|3176_ , \new_Sorter100|3177_ , \new_Sorter100|3178_ ,
    \new_Sorter100|3179_ , \new_Sorter100|3180_ , \new_Sorter100|3181_ ,
    \new_Sorter100|3182_ , \new_Sorter100|3183_ , \new_Sorter100|3184_ ,
    \new_Sorter100|3185_ , \new_Sorter100|3186_ , \new_Sorter100|3187_ ,
    \new_Sorter100|3188_ , \new_Sorter100|3189_ , \new_Sorter100|3190_ ,
    \new_Sorter100|3191_ , \new_Sorter100|3192_ , \new_Sorter100|3193_ ,
    \new_Sorter100|3194_ , \new_Sorter100|3195_ , \new_Sorter100|3196_ ,
    \new_Sorter100|3197_ , \new_Sorter100|3198_ , \new_Sorter100|3200_ ,
    \new_Sorter100|3201_ , \new_Sorter100|3202_ , \new_Sorter100|3203_ ,
    \new_Sorter100|3204_ , \new_Sorter100|3205_ , \new_Sorter100|3206_ ,
    \new_Sorter100|3207_ , \new_Sorter100|3208_ , \new_Sorter100|3209_ ,
    \new_Sorter100|3210_ , \new_Sorter100|3211_ , \new_Sorter100|3212_ ,
    \new_Sorter100|3213_ , \new_Sorter100|3214_ , \new_Sorter100|3215_ ,
    \new_Sorter100|3216_ , \new_Sorter100|3217_ , \new_Sorter100|3218_ ,
    \new_Sorter100|3219_ , \new_Sorter100|3220_ , \new_Sorter100|3221_ ,
    \new_Sorter100|3222_ , \new_Sorter100|3223_ , \new_Sorter100|3224_ ,
    \new_Sorter100|3225_ , \new_Sorter100|3226_ , \new_Sorter100|3227_ ,
    \new_Sorter100|3228_ , \new_Sorter100|3229_ , \new_Sorter100|3230_ ,
    \new_Sorter100|3231_ , \new_Sorter100|3232_ , \new_Sorter100|3233_ ,
    \new_Sorter100|3234_ , \new_Sorter100|3235_ , \new_Sorter100|3236_ ,
    \new_Sorter100|3237_ , \new_Sorter100|3238_ , \new_Sorter100|3239_ ,
    \new_Sorter100|3240_ , \new_Sorter100|3241_ , \new_Sorter100|3242_ ,
    \new_Sorter100|3243_ , \new_Sorter100|3244_ , \new_Sorter100|3245_ ,
    \new_Sorter100|3246_ , \new_Sorter100|3247_ , \new_Sorter100|3248_ ,
    \new_Sorter100|3249_ , \new_Sorter100|3250_ , \new_Sorter100|3251_ ,
    \new_Sorter100|3252_ , \new_Sorter100|3253_ , \new_Sorter100|3254_ ,
    \new_Sorter100|3255_ , \new_Sorter100|3256_ , \new_Sorter100|3257_ ,
    \new_Sorter100|3258_ , \new_Sorter100|3259_ , \new_Sorter100|3260_ ,
    \new_Sorter100|3261_ , \new_Sorter100|3262_ , \new_Sorter100|3263_ ,
    \new_Sorter100|3264_ , \new_Sorter100|3265_ , \new_Sorter100|3266_ ,
    \new_Sorter100|3267_ , \new_Sorter100|3268_ , \new_Sorter100|3269_ ,
    \new_Sorter100|3270_ , \new_Sorter100|3271_ , \new_Sorter100|3272_ ,
    \new_Sorter100|3273_ , \new_Sorter100|3274_ , \new_Sorter100|3275_ ,
    \new_Sorter100|3276_ , \new_Sorter100|3277_ , \new_Sorter100|3278_ ,
    \new_Sorter100|3279_ , \new_Sorter100|3280_ , \new_Sorter100|3281_ ,
    \new_Sorter100|3282_ , \new_Sorter100|3283_ , \new_Sorter100|3284_ ,
    \new_Sorter100|3285_ , \new_Sorter100|3286_ , \new_Sorter100|3287_ ,
    \new_Sorter100|3288_ , \new_Sorter100|3289_ , \new_Sorter100|3290_ ,
    \new_Sorter100|3291_ , \new_Sorter100|3292_ , \new_Sorter100|3293_ ,
    \new_Sorter100|3294_ , \new_Sorter100|3295_ , \new_Sorter100|3296_ ,
    \new_Sorter100|3297_ , \new_Sorter100|3298_ , \new_Sorter100|3299_ ,
    \new_Sorter100|3300_ , \new_Sorter100|3399_ , \new_Sorter100|3301_ ,
    \new_Sorter100|3302_ , \new_Sorter100|3303_ , \new_Sorter100|3304_ ,
    \new_Sorter100|3305_ , \new_Sorter100|3306_ , \new_Sorter100|3307_ ,
    \new_Sorter100|3308_ , \new_Sorter100|3309_ , \new_Sorter100|3310_ ,
    \new_Sorter100|3311_ , \new_Sorter100|3312_ , \new_Sorter100|3313_ ,
    \new_Sorter100|3314_ , \new_Sorter100|3315_ , \new_Sorter100|3316_ ,
    \new_Sorter100|3317_ , \new_Sorter100|3318_ , \new_Sorter100|3319_ ,
    \new_Sorter100|3320_ , \new_Sorter100|3321_ , \new_Sorter100|3322_ ,
    \new_Sorter100|3323_ , \new_Sorter100|3324_ , \new_Sorter100|3325_ ,
    \new_Sorter100|3326_ , \new_Sorter100|3327_ , \new_Sorter100|3328_ ,
    \new_Sorter100|3329_ , \new_Sorter100|3330_ , \new_Sorter100|3331_ ,
    \new_Sorter100|3332_ , \new_Sorter100|3333_ , \new_Sorter100|3334_ ,
    \new_Sorter100|3335_ , \new_Sorter100|3336_ , \new_Sorter100|3337_ ,
    \new_Sorter100|3338_ , \new_Sorter100|3339_ , \new_Sorter100|3340_ ,
    \new_Sorter100|3341_ , \new_Sorter100|3342_ , \new_Sorter100|3343_ ,
    \new_Sorter100|3344_ , \new_Sorter100|3345_ , \new_Sorter100|3346_ ,
    \new_Sorter100|3347_ , \new_Sorter100|3348_ , \new_Sorter100|3349_ ,
    \new_Sorter100|3350_ , \new_Sorter100|3351_ , \new_Sorter100|3352_ ,
    \new_Sorter100|3353_ , \new_Sorter100|3354_ , \new_Sorter100|3355_ ,
    \new_Sorter100|3356_ , \new_Sorter100|3357_ , \new_Sorter100|3358_ ,
    \new_Sorter100|3359_ , \new_Sorter100|3360_ , \new_Sorter100|3361_ ,
    \new_Sorter100|3362_ , \new_Sorter100|3363_ , \new_Sorter100|3364_ ,
    \new_Sorter100|3365_ , \new_Sorter100|3366_ , \new_Sorter100|3367_ ,
    \new_Sorter100|3368_ , \new_Sorter100|3369_ , \new_Sorter100|3370_ ,
    \new_Sorter100|3371_ , \new_Sorter100|3372_ , \new_Sorter100|3373_ ,
    \new_Sorter100|3374_ , \new_Sorter100|3375_ , \new_Sorter100|3376_ ,
    \new_Sorter100|3377_ , \new_Sorter100|3378_ , \new_Sorter100|3379_ ,
    \new_Sorter100|3380_ , \new_Sorter100|3381_ , \new_Sorter100|3382_ ,
    \new_Sorter100|3383_ , \new_Sorter100|3384_ , \new_Sorter100|3385_ ,
    \new_Sorter100|3386_ , \new_Sorter100|3387_ , \new_Sorter100|3388_ ,
    \new_Sorter100|3389_ , \new_Sorter100|3390_ , \new_Sorter100|3391_ ,
    \new_Sorter100|3392_ , \new_Sorter100|3393_ , \new_Sorter100|3394_ ,
    \new_Sorter100|3395_ , \new_Sorter100|3396_ , \new_Sorter100|3397_ ,
    \new_Sorter100|3398_ , \new_Sorter100|3400_ , \new_Sorter100|3401_ ,
    \new_Sorter100|3402_ , \new_Sorter100|3403_ , \new_Sorter100|3404_ ,
    \new_Sorter100|3405_ , \new_Sorter100|3406_ , \new_Sorter100|3407_ ,
    \new_Sorter100|3408_ , \new_Sorter100|3409_ , \new_Sorter100|3410_ ,
    \new_Sorter100|3411_ , \new_Sorter100|3412_ , \new_Sorter100|3413_ ,
    \new_Sorter100|3414_ , \new_Sorter100|3415_ , \new_Sorter100|3416_ ,
    \new_Sorter100|3417_ , \new_Sorter100|3418_ , \new_Sorter100|3419_ ,
    \new_Sorter100|3420_ , \new_Sorter100|3421_ , \new_Sorter100|3422_ ,
    \new_Sorter100|3423_ , \new_Sorter100|3424_ , \new_Sorter100|3425_ ,
    \new_Sorter100|3426_ , \new_Sorter100|3427_ , \new_Sorter100|3428_ ,
    \new_Sorter100|3429_ , \new_Sorter100|3430_ , \new_Sorter100|3431_ ,
    \new_Sorter100|3432_ , \new_Sorter100|3433_ , \new_Sorter100|3434_ ,
    \new_Sorter100|3435_ , \new_Sorter100|3436_ , \new_Sorter100|3437_ ,
    \new_Sorter100|3438_ , \new_Sorter100|3439_ , \new_Sorter100|3440_ ,
    \new_Sorter100|3441_ , \new_Sorter100|3442_ , \new_Sorter100|3443_ ,
    \new_Sorter100|3444_ , \new_Sorter100|3445_ , \new_Sorter100|3446_ ,
    \new_Sorter100|3447_ , \new_Sorter100|3448_ , \new_Sorter100|3449_ ,
    \new_Sorter100|3450_ , \new_Sorter100|3451_ , \new_Sorter100|3452_ ,
    \new_Sorter100|3453_ , \new_Sorter100|3454_ , \new_Sorter100|3455_ ,
    \new_Sorter100|3456_ , \new_Sorter100|3457_ , \new_Sorter100|3458_ ,
    \new_Sorter100|3459_ , \new_Sorter100|3460_ , \new_Sorter100|3461_ ,
    \new_Sorter100|3462_ , \new_Sorter100|3463_ , \new_Sorter100|3464_ ,
    \new_Sorter100|3465_ , \new_Sorter100|3466_ , \new_Sorter100|3467_ ,
    \new_Sorter100|3468_ , \new_Sorter100|3469_ , \new_Sorter100|3470_ ,
    \new_Sorter100|3471_ , \new_Sorter100|3472_ , \new_Sorter100|3473_ ,
    \new_Sorter100|3474_ , \new_Sorter100|3475_ , \new_Sorter100|3476_ ,
    \new_Sorter100|3477_ , \new_Sorter100|3478_ , \new_Sorter100|3479_ ,
    \new_Sorter100|3480_ , \new_Sorter100|3481_ , \new_Sorter100|3482_ ,
    \new_Sorter100|3483_ , \new_Sorter100|3484_ , \new_Sorter100|3485_ ,
    \new_Sorter100|3486_ , \new_Sorter100|3487_ , \new_Sorter100|3488_ ,
    \new_Sorter100|3489_ , \new_Sorter100|3490_ , \new_Sorter100|3491_ ,
    \new_Sorter100|3492_ , \new_Sorter100|3493_ , \new_Sorter100|3494_ ,
    \new_Sorter100|3495_ , \new_Sorter100|3496_ , \new_Sorter100|3497_ ,
    \new_Sorter100|3498_ , \new_Sorter100|3499_ , \new_Sorter100|3500_ ,
    \new_Sorter100|3599_ , \new_Sorter100|3501_ , \new_Sorter100|3502_ ,
    \new_Sorter100|3503_ , \new_Sorter100|3504_ , \new_Sorter100|3505_ ,
    \new_Sorter100|3506_ , \new_Sorter100|3507_ , \new_Sorter100|3508_ ,
    \new_Sorter100|3509_ , \new_Sorter100|3510_ , \new_Sorter100|3511_ ,
    \new_Sorter100|3512_ , \new_Sorter100|3513_ , \new_Sorter100|3514_ ,
    \new_Sorter100|3515_ , \new_Sorter100|3516_ , \new_Sorter100|3517_ ,
    \new_Sorter100|3518_ , \new_Sorter100|3519_ , \new_Sorter100|3520_ ,
    \new_Sorter100|3521_ , \new_Sorter100|3522_ , \new_Sorter100|3523_ ,
    \new_Sorter100|3524_ , \new_Sorter100|3525_ , \new_Sorter100|3526_ ,
    \new_Sorter100|3527_ , \new_Sorter100|3528_ , \new_Sorter100|3529_ ,
    \new_Sorter100|3530_ , \new_Sorter100|3531_ , \new_Sorter100|3532_ ,
    \new_Sorter100|3533_ , \new_Sorter100|3534_ , \new_Sorter100|3535_ ,
    \new_Sorter100|3536_ , \new_Sorter100|3537_ , \new_Sorter100|3538_ ,
    \new_Sorter100|3539_ , \new_Sorter100|3540_ , \new_Sorter100|3541_ ,
    \new_Sorter100|3542_ , \new_Sorter100|3543_ , \new_Sorter100|3544_ ,
    \new_Sorter100|3545_ , \new_Sorter100|3546_ , \new_Sorter100|3547_ ,
    \new_Sorter100|3548_ , \new_Sorter100|3549_ , \new_Sorter100|3550_ ,
    \new_Sorter100|3551_ , \new_Sorter100|3552_ , \new_Sorter100|3553_ ,
    \new_Sorter100|3554_ , \new_Sorter100|3555_ , \new_Sorter100|3556_ ,
    \new_Sorter100|3557_ , \new_Sorter100|3558_ , \new_Sorter100|3559_ ,
    \new_Sorter100|3560_ , \new_Sorter100|3561_ , \new_Sorter100|3562_ ,
    \new_Sorter100|3563_ , \new_Sorter100|3564_ , \new_Sorter100|3565_ ,
    \new_Sorter100|3566_ , \new_Sorter100|3567_ , \new_Sorter100|3568_ ,
    \new_Sorter100|3569_ , \new_Sorter100|3570_ , \new_Sorter100|3571_ ,
    \new_Sorter100|3572_ , \new_Sorter100|3573_ , \new_Sorter100|3574_ ,
    \new_Sorter100|3575_ , \new_Sorter100|3576_ , \new_Sorter100|3577_ ,
    \new_Sorter100|3578_ , \new_Sorter100|3579_ , \new_Sorter100|3580_ ,
    \new_Sorter100|3581_ , \new_Sorter100|3582_ , \new_Sorter100|3583_ ,
    \new_Sorter100|3584_ , \new_Sorter100|3585_ , \new_Sorter100|3586_ ,
    \new_Sorter100|3587_ , \new_Sorter100|3588_ , \new_Sorter100|3589_ ,
    \new_Sorter100|3590_ , \new_Sorter100|3591_ , \new_Sorter100|3592_ ,
    \new_Sorter100|3593_ , \new_Sorter100|3594_ , \new_Sorter100|3595_ ,
    \new_Sorter100|3596_ , \new_Sorter100|3597_ , \new_Sorter100|3598_ ,
    \new_Sorter100|3600_ , \new_Sorter100|3601_ , \new_Sorter100|3602_ ,
    \new_Sorter100|3603_ , \new_Sorter100|3604_ , \new_Sorter100|3605_ ,
    \new_Sorter100|3606_ , \new_Sorter100|3607_ , \new_Sorter100|3608_ ,
    \new_Sorter100|3609_ , \new_Sorter100|3610_ , \new_Sorter100|3611_ ,
    \new_Sorter100|3612_ , \new_Sorter100|3613_ , \new_Sorter100|3614_ ,
    \new_Sorter100|3615_ , \new_Sorter100|3616_ , \new_Sorter100|3617_ ,
    \new_Sorter100|3618_ , \new_Sorter100|3619_ , \new_Sorter100|3620_ ,
    \new_Sorter100|3621_ , \new_Sorter100|3622_ , \new_Sorter100|3623_ ,
    \new_Sorter100|3624_ , \new_Sorter100|3625_ , \new_Sorter100|3626_ ,
    \new_Sorter100|3627_ , \new_Sorter100|3628_ , \new_Sorter100|3629_ ,
    \new_Sorter100|3630_ , \new_Sorter100|3631_ , \new_Sorter100|3632_ ,
    \new_Sorter100|3633_ , \new_Sorter100|3634_ , \new_Sorter100|3635_ ,
    \new_Sorter100|3636_ , \new_Sorter100|3637_ , \new_Sorter100|3638_ ,
    \new_Sorter100|3639_ , \new_Sorter100|3640_ , \new_Sorter100|3641_ ,
    \new_Sorter100|3642_ , \new_Sorter100|3643_ , \new_Sorter100|3644_ ,
    \new_Sorter100|3645_ , \new_Sorter100|3646_ , \new_Sorter100|3647_ ,
    \new_Sorter100|3648_ , \new_Sorter100|3649_ , \new_Sorter100|3650_ ,
    \new_Sorter100|3651_ , \new_Sorter100|3652_ , \new_Sorter100|3653_ ,
    \new_Sorter100|3654_ , \new_Sorter100|3655_ , \new_Sorter100|3656_ ,
    \new_Sorter100|3657_ , \new_Sorter100|3658_ , \new_Sorter100|3659_ ,
    \new_Sorter100|3660_ , \new_Sorter100|3661_ , \new_Sorter100|3662_ ,
    \new_Sorter100|3663_ , \new_Sorter100|3664_ , \new_Sorter100|3665_ ,
    \new_Sorter100|3666_ , \new_Sorter100|3667_ , \new_Sorter100|3668_ ,
    \new_Sorter100|3669_ , \new_Sorter100|3670_ , \new_Sorter100|3671_ ,
    \new_Sorter100|3672_ , \new_Sorter100|3673_ , \new_Sorter100|3674_ ,
    \new_Sorter100|3675_ , \new_Sorter100|3676_ , \new_Sorter100|3677_ ,
    \new_Sorter100|3678_ , \new_Sorter100|3679_ , \new_Sorter100|3680_ ,
    \new_Sorter100|3681_ , \new_Sorter100|3682_ , \new_Sorter100|3683_ ,
    \new_Sorter100|3684_ , \new_Sorter100|3685_ , \new_Sorter100|3686_ ,
    \new_Sorter100|3687_ , \new_Sorter100|3688_ , \new_Sorter100|3689_ ,
    \new_Sorter100|3690_ , \new_Sorter100|3691_ , \new_Sorter100|3692_ ,
    \new_Sorter100|3693_ , \new_Sorter100|3694_ , \new_Sorter100|3695_ ,
    \new_Sorter100|3696_ , \new_Sorter100|3697_ , \new_Sorter100|3698_ ,
    \new_Sorter100|3699_ , \new_Sorter100|3700_ , \new_Sorter100|3799_ ,
    \new_Sorter100|3701_ , \new_Sorter100|3702_ , \new_Sorter100|3703_ ,
    \new_Sorter100|3704_ , \new_Sorter100|3705_ , \new_Sorter100|3706_ ,
    \new_Sorter100|3707_ , \new_Sorter100|3708_ , \new_Sorter100|3709_ ,
    \new_Sorter100|3710_ , \new_Sorter100|3711_ , \new_Sorter100|3712_ ,
    \new_Sorter100|3713_ , \new_Sorter100|3714_ , \new_Sorter100|3715_ ,
    \new_Sorter100|3716_ , \new_Sorter100|3717_ , \new_Sorter100|3718_ ,
    \new_Sorter100|3719_ , \new_Sorter100|3720_ , \new_Sorter100|3721_ ,
    \new_Sorter100|3722_ , \new_Sorter100|3723_ , \new_Sorter100|3724_ ,
    \new_Sorter100|3725_ , \new_Sorter100|3726_ , \new_Sorter100|3727_ ,
    \new_Sorter100|3728_ , \new_Sorter100|3729_ , \new_Sorter100|3730_ ,
    \new_Sorter100|3731_ , \new_Sorter100|3732_ , \new_Sorter100|3733_ ,
    \new_Sorter100|3734_ , \new_Sorter100|3735_ , \new_Sorter100|3736_ ,
    \new_Sorter100|3737_ , \new_Sorter100|3738_ , \new_Sorter100|3739_ ,
    \new_Sorter100|3740_ , \new_Sorter100|3741_ , \new_Sorter100|3742_ ,
    \new_Sorter100|3743_ , \new_Sorter100|3744_ , \new_Sorter100|3745_ ,
    \new_Sorter100|3746_ , \new_Sorter100|3747_ , \new_Sorter100|3748_ ,
    \new_Sorter100|3749_ , \new_Sorter100|3750_ , \new_Sorter100|3751_ ,
    \new_Sorter100|3752_ , \new_Sorter100|3753_ , \new_Sorter100|3754_ ,
    \new_Sorter100|3755_ , \new_Sorter100|3756_ , \new_Sorter100|3757_ ,
    \new_Sorter100|3758_ , \new_Sorter100|3759_ , \new_Sorter100|3760_ ,
    \new_Sorter100|3761_ , \new_Sorter100|3762_ , \new_Sorter100|3763_ ,
    \new_Sorter100|3764_ , \new_Sorter100|3765_ , \new_Sorter100|3766_ ,
    \new_Sorter100|3767_ , \new_Sorter100|3768_ , \new_Sorter100|3769_ ,
    \new_Sorter100|3770_ , \new_Sorter100|3771_ , \new_Sorter100|3772_ ,
    \new_Sorter100|3773_ , \new_Sorter100|3774_ , \new_Sorter100|3775_ ,
    \new_Sorter100|3776_ , \new_Sorter100|3777_ , \new_Sorter100|3778_ ,
    \new_Sorter100|3779_ , \new_Sorter100|3780_ , \new_Sorter100|3781_ ,
    \new_Sorter100|3782_ , \new_Sorter100|3783_ , \new_Sorter100|3784_ ,
    \new_Sorter100|3785_ , \new_Sorter100|3786_ , \new_Sorter100|3787_ ,
    \new_Sorter100|3788_ , \new_Sorter100|3789_ , \new_Sorter100|3790_ ,
    \new_Sorter100|3791_ , \new_Sorter100|3792_ , \new_Sorter100|3793_ ,
    \new_Sorter100|3794_ , \new_Sorter100|3795_ , \new_Sorter100|3796_ ,
    \new_Sorter100|3797_ , \new_Sorter100|3798_ , \new_Sorter100|3800_ ,
    \new_Sorter100|3801_ , \new_Sorter100|3802_ , \new_Sorter100|3803_ ,
    \new_Sorter100|3804_ , \new_Sorter100|3805_ , \new_Sorter100|3806_ ,
    \new_Sorter100|3807_ , \new_Sorter100|3808_ , \new_Sorter100|3809_ ,
    \new_Sorter100|3810_ , \new_Sorter100|3811_ , \new_Sorter100|3812_ ,
    \new_Sorter100|3813_ , \new_Sorter100|3814_ , \new_Sorter100|3815_ ,
    \new_Sorter100|3816_ , \new_Sorter100|3817_ , \new_Sorter100|3818_ ,
    \new_Sorter100|3819_ , \new_Sorter100|3820_ , \new_Sorter100|3821_ ,
    \new_Sorter100|3822_ , \new_Sorter100|3823_ , \new_Sorter100|3824_ ,
    \new_Sorter100|3825_ , \new_Sorter100|3826_ , \new_Sorter100|3827_ ,
    \new_Sorter100|3828_ , \new_Sorter100|3829_ , \new_Sorter100|3830_ ,
    \new_Sorter100|3831_ , \new_Sorter100|3832_ , \new_Sorter100|3833_ ,
    \new_Sorter100|3834_ , \new_Sorter100|3835_ , \new_Sorter100|3836_ ,
    \new_Sorter100|3837_ , \new_Sorter100|3838_ , \new_Sorter100|3839_ ,
    \new_Sorter100|3840_ , \new_Sorter100|3841_ , \new_Sorter100|3842_ ,
    \new_Sorter100|3843_ , \new_Sorter100|3844_ , \new_Sorter100|3845_ ,
    \new_Sorter100|3846_ , \new_Sorter100|3847_ , \new_Sorter100|3848_ ,
    \new_Sorter100|3849_ , \new_Sorter100|3850_ , \new_Sorter100|3851_ ,
    \new_Sorter100|3852_ , \new_Sorter100|3853_ , \new_Sorter100|3854_ ,
    \new_Sorter100|3855_ , \new_Sorter100|3856_ , \new_Sorter100|3857_ ,
    \new_Sorter100|3858_ , \new_Sorter100|3859_ , \new_Sorter100|3860_ ,
    \new_Sorter100|3861_ , \new_Sorter100|3862_ , \new_Sorter100|3863_ ,
    \new_Sorter100|3864_ , \new_Sorter100|3865_ , \new_Sorter100|3866_ ,
    \new_Sorter100|3867_ , \new_Sorter100|3868_ , \new_Sorter100|3869_ ,
    \new_Sorter100|3870_ , \new_Sorter100|3871_ , \new_Sorter100|3872_ ,
    \new_Sorter100|3873_ , \new_Sorter100|3874_ , \new_Sorter100|3875_ ,
    \new_Sorter100|3876_ , \new_Sorter100|3877_ , \new_Sorter100|3878_ ,
    \new_Sorter100|3879_ , \new_Sorter100|3880_ , \new_Sorter100|3881_ ,
    \new_Sorter100|3882_ , \new_Sorter100|3883_ , \new_Sorter100|3884_ ,
    \new_Sorter100|3885_ , \new_Sorter100|3886_ , \new_Sorter100|3887_ ,
    \new_Sorter100|3888_ , \new_Sorter100|3889_ , \new_Sorter100|3890_ ,
    \new_Sorter100|3891_ , \new_Sorter100|3892_ , \new_Sorter100|3893_ ,
    \new_Sorter100|3894_ , \new_Sorter100|3895_ , \new_Sorter100|3896_ ,
    \new_Sorter100|3897_ , \new_Sorter100|3898_ , \new_Sorter100|3899_ ,
    \new_Sorter100|3900_ , \new_Sorter100|3999_ , \new_Sorter100|3901_ ,
    \new_Sorter100|3902_ , \new_Sorter100|3903_ , \new_Sorter100|3904_ ,
    \new_Sorter100|3905_ , \new_Sorter100|3906_ , \new_Sorter100|3907_ ,
    \new_Sorter100|3908_ , \new_Sorter100|3909_ , \new_Sorter100|3910_ ,
    \new_Sorter100|3911_ , \new_Sorter100|3912_ , \new_Sorter100|3913_ ,
    \new_Sorter100|3914_ , \new_Sorter100|3915_ , \new_Sorter100|3916_ ,
    \new_Sorter100|3917_ , \new_Sorter100|3918_ , \new_Sorter100|3919_ ,
    \new_Sorter100|3920_ , \new_Sorter100|3921_ , \new_Sorter100|3922_ ,
    \new_Sorter100|3923_ , \new_Sorter100|3924_ , \new_Sorter100|3925_ ,
    \new_Sorter100|3926_ , \new_Sorter100|3927_ , \new_Sorter100|3928_ ,
    \new_Sorter100|3929_ , \new_Sorter100|3930_ , \new_Sorter100|3931_ ,
    \new_Sorter100|3932_ , \new_Sorter100|3933_ , \new_Sorter100|3934_ ,
    \new_Sorter100|3935_ , \new_Sorter100|3936_ , \new_Sorter100|3937_ ,
    \new_Sorter100|3938_ , \new_Sorter100|3939_ , \new_Sorter100|3940_ ,
    \new_Sorter100|3941_ , \new_Sorter100|3942_ , \new_Sorter100|3943_ ,
    \new_Sorter100|3944_ , \new_Sorter100|3945_ , \new_Sorter100|3946_ ,
    \new_Sorter100|3947_ , \new_Sorter100|3948_ , \new_Sorter100|3949_ ,
    \new_Sorter100|3950_ , \new_Sorter100|3951_ , \new_Sorter100|3952_ ,
    \new_Sorter100|3953_ , \new_Sorter100|3954_ , \new_Sorter100|3955_ ,
    \new_Sorter100|3956_ , \new_Sorter100|3957_ , \new_Sorter100|3958_ ,
    \new_Sorter100|3959_ , \new_Sorter100|3960_ , \new_Sorter100|3961_ ,
    \new_Sorter100|3962_ , \new_Sorter100|3963_ , \new_Sorter100|3964_ ,
    \new_Sorter100|3965_ , \new_Sorter100|3966_ , \new_Sorter100|3967_ ,
    \new_Sorter100|3968_ , \new_Sorter100|3969_ , \new_Sorter100|3970_ ,
    \new_Sorter100|3971_ , \new_Sorter100|3972_ , \new_Sorter100|3973_ ,
    \new_Sorter100|3974_ , \new_Sorter100|3975_ , \new_Sorter100|3976_ ,
    \new_Sorter100|3977_ , \new_Sorter100|3978_ , \new_Sorter100|3979_ ,
    \new_Sorter100|3980_ , \new_Sorter100|3981_ , \new_Sorter100|3982_ ,
    \new_Sorter100|3983_ , \new_Sorter100|3984_ , \new_Sorter100|3985_ ,
    \new_Sorter100|3986_ , \new_Sorter100|3987_ , \new_Sorter100|3988_ ,
    \new_Sorter100|3989_ , \new_Sorter100|3990_ , \new_Sorter100|3991_ ,
    \new_Sorter100|3992_ , \new_Sorter100|3993_ , \new_Sorter100|3994_ ,
    \new_Sorter100|3995_ , \new_Sorter100|3996_ , \new_Sorter100|3997_ ,
    \new_Sorter100|3998_ , \new_Sorter100|4000_ , \new_Sorter100|4001_ ,
    \new_Sorter100|4002_ , \new_Sorter100|4003_ , \new_Sorter100|4004_ ,
    \new_Sorter100|4005_ , \new_Sorter100|4006_ , \new_Sorter100|4007_ ,
    \new_Sorter100|4008_ , \new_Sorter100|4009_ , \new_Sorter100|4010_ ,
    \new_Sorter100|4011_ , \new_Sorter100|4012_ , \new_Sorter100|4013_ ,
    \new_Sorter100|4014_ , \new_Sorter100|4015_ , \new_Sorter100|4016_ ,
    \new_Sorter100|4017_ , \new_Sorter100|4018_ , \new_Sorter100|4019_ ,
    \new_Sorter100|4020_ , \new_Sorter100|4021_ , \new_Sorter100|4022_ ,
    \new_Sorter100|4023_ , \new_Sorter100|4024_ , \new_Sorter100|4025_ ,
    \new_Sorter100|4026_ , \new_Sorter100|4027_ , \new_Sorter100|4028_ ,
    \new_Sorter100|4029_ , \new_Sorter100|4030_ , \new_Sorter100|4031_ ,
    \new_Sorter100|4032_ , \new_Sorter100|4033_ , \new_Sorter100|4034_ ,
    \new_Sorter100|4035_ , \new_Sorter100|4036_ , \new_Sorter100|4037_ ,
    \new_Sorter100|4038_ , \new_Sorter100|4039_ , \new_Sorter100|4040_ ,
    \new_Sorter100|4041_ , \new_Sorter100|4042_ , \new_Sorter100|4043_ ,
    \new_Sorter100|4044_ , \new_Sorter100|4045_ , \new_Sorter100|4046_ ,
    \new_Sorter100|4047_ , \new_Sorter100|4048_ , \new_Sorter100|4049_ ,
    \new_Sorter100|4050_ , \new_Sorter100|4051_ , \new_Sorter100|4052_ ,
    \new_Sorter100|4053_ , \new_Sorter100|4054_ , \new_Sorter100|4055_ ,
    \new_Sorter100|4056_ , \new_Sorter100|4057_ , \new_Sorter100|4058_ ,
    \new_Sorter100|4059_ , \new_Sorter100|4060_ , \new_Sorter100|4061_ ,
    \new_Sorter100|4062_ , \new_Sorter100|4063_ , \new_Sorter100|4064_ ,
    \new_Sorter100|4065_ , \new_Sorter100|4066_ , \new_Sorter100|4067_ ,
    \new_Sorter100|4068_ , \new_Sorter100|4069_ , \new_Sorter100|4070_ ,
    \new_Sorter100|4071_ , \new_Sorter100|4072_ , \new_Sorter100|4073_ ,
    \new_Sorter100|4074_ , \new_Sorter100|4075_ , \new_Sorter100|4076_ ,
    \new_Sorter100|4077_ , \new_Sorter100|4078_ , \new_Sorter100|4079_ ,
    \new_Sorter100|4080_ , \new_Sorter100|4081_ , \new_Sorter100|4082_ ,
    \new_Sorter100|4083_ , \new_Sorter100|4084_ , \new_Sorter100|4085_ ,
    \new_Sorter100|4086_ , \new_Sorter100|4087_ , \new_Sorter100|4088_ ,
    \new_Sorter100|4089_ , \new_Sorter100|4090_ , \new_Sorter100|4091_ ,
    \new_Sorter100|4092_ , \new_Sorter100|4093_ , \new_Sorter100|4094_ ,
    \new_Sorter100|4095_ , \new_Sorter100|4096_ , \new_Sorter100|4097_ ,
    \new_Sorter100|4098_ , \new_Sorter100|4099_ , \new_Sorter100|4100_ ,
    \new_Sorter100|4199_ , \new_Sorter100|4101_ , \new_Sorter100|4102_ ,
    \new_Sorter100|4103_ , \new_Sorter100|4104_ , \new_Sorter100|4105_ ,
    \new_Sorter100|4106_ , \new_Sorter100|4107_ , \new_Sorter100|4108_ ,
    \new_Sorter100|4109_ , \new_Sorter100|4110_ , \new_Sorter100|4111_ ,
    \new_Sorter100|4112_ , \new_Sorter100|4113_ , \new_Sorter100|4114_ ,
    \new_Sorter100|4115_ , \new_Sorter100|4116_ , \new_Sorter100|4117_ ,
    \new_Sorter100|4118_ , \new_Sorter100|4119_ , \new_Sorter100|4120_ ,
    \new_Sorter100|4121_ , \new_Sorter100|4122_ , \new_Sorter100|4123_ ,
    \new_Sorter100|4124_ , \new_Sorter100|4125_ , \new_Sorter100|4126_ ,
    \new_Sorter100|4127_ , \new_Sorter100|4128_ , \new_Sorter100|4129_ ,
    \new_Sorter100|4130_ , \new_Sorter100|4131_ , \new_Sorter100|4132_ ,
    \new_Sorter100|4133_ , \new_Sorter100|4134_ , \new_Sorter100|4135_ ,
    \new_Sorter100|4136_ , \new_Sorter100|4137_ , \new_Sorter100|4138_ ,
    \new_Sorter100|4139_ , \new_Sorter100|4140_ , \new_Sorter100|4141_ ,
    \new_Sorter100|4142_ , \new_Sorter100|4143_ , \new_Sorter100|4144_ ,
    \new_Sorter100|4145_ , \new_Sorter100|4146_ , \new_Sorter100|4147_ ,
    \new_Sorter100|4148_ , \new_Sorter100|4149_ , \new_Sorter100|4150_ ,
    \new_Sorter100|4151_ , \new_Sorter100|4152_ , \new_Sorter100|4153_ ,
    \new_Sorter100|4154_ , \new_Sorter100|4155_ , \new_Sorter100|4156_ ,
    \new_Sorter100|4157_ , \new_Sorter100|4158_ , \new_Sorter100|4159_ ,
    \new_Sorter100|4160_ , \new_Sorter100|4161_ , \new_Sorter100|4162_ ,
    \new_Sorter100|4163_ , \new_Sorter100|4164_ , \new_Sorter100|4165_ ,
    \new_Sorter100|4166_ , \new_Sorter100|4167_ , \new_Sorter100|4168_ ,
    \new_Sorter100|4169_ , \new_Sorter100|4170_ , \new_Sorter100|4171_ ,
    \new_Sorter100|4172_ , \new_Sorter100|4173_ , \new_Sorter100|4174_ ,
    \new_Sorter100|4175_ , \new_Sorter100|4176_ , \new_Sorter100|4177_ ,
    \new_Sorter100|4178_ , \new_Sorter100|4179_ , \new_Sorter100|4180_ ,
    \new_Sorter100|4181_ , \new_Sorter100|4182_ , \new_Sorter100|4183_ ,
    \new_Sorter100|4184_ , \new_Sorter100|4185_ , \new_Sorter100|4186_ ,
    \new_Sorter100|4187_ , \new_Sorter100|4188_ , \new_Sorter100|4189_ ,
    \new_Sorter100|4190_ , \new_Sorter100|4191_ , \new_Sorter100|4192_ ,
    \new_Sorter100|4193_ , \new_Sorter100|4194_ , \new_Sorter100|4195_ ,
    \new_Sorter100|4196_ , \new_Sorter100|4197_ , \new_Sorter100|4198_ ,
    \new_Sorter100|4200_ , \new_Sorter100|4201_ , \new_Sorter100|4202_ ,
    \new_Sorter100|4203_ , \new_Sorter100|4204_ , \new_Sorter100|4205_ ,
    \new_Sorter100|4206_ , \new_Sorter100|4207_ , \new_Sorter100|4208_ ,
    \new_Sorter100|4209_ , \new_Sorter100|4210_ , \new_Sorter100|4211_ ,
    \new_Sorter100|4212_ , \new_Sorter100|4213_ , \new_Sorter100|4214_ ,
    \new_Sorter100|4215_ , \new_Sorter100|4216_ , \new_Sorter100|4217_ ,
    \new_Sorter100|4218_ , \new_Sorter100|4219_ , \new_Sorter100|4220_ ,
    \new_Sorter100|4221_ , \new_Sorter100|4222_ , \new_Sorter100|4223_ ,
    \new_Sorter100|4224_ , \new_Sorter100|4225_ , \new_Sorter100|4226_ ,
    \new_Sorter100|4227_ , \new_Sorter100|4228_ , \new_Sorter100|4229_ ,
    \new_Sorter100|4230_ , \new_Sorter100|4231_ , \new_Sorter100|4232_ ,
    \new_Sorter100|4233_ , \new_Sorter100|4234_ , \new_Sorter100|4235_ ,
    \new_Sorter100|4236_ , \new_Sorter100|4237_ , \new_Sorter100|4238_ ,
    \new_Sorter100|4239_ , \new_Sorter100|4240_ , \new_Sorter100|4241_ ,
    \new_Sorter100|4242_ , \new_Sorter100|4243_ , \new_Sorter100|4244_ ,
    \new_Sorter100|4245_ , \new_Sorter100|4246_ , \new_Sorter100|4247_ ,
    \new_Sorter100|4248_ , \new_Sorter100|4249_ , \new_Sorter100|4250_ ,
    \new_Sorter100|4251_ , \new_Sorter100|4252_ , \new_Sorter100|4253_ ,
    \new_Sorter100|4254_ , \new_Sorter100|4255_ , \new_Sorter100|4256_ ,
    \new_Sorter100|4257_ , \new_Sorter100|4258_ , \new_Sorter100|4259_ ,
    \new_Sorter100|4260_ , \new_Sorter100|4261_ , \new_Sorter100|4262_ ,
    \new_Sorter100|4263_ , \new_Sorter100|4264_ , \new_Sorter100|4265_ ,
    \new_Sorter100|4266_ , \new_Sorter100|4267_ , \new_Sorter100|4268_ ,
    \new_Sorter100|4269_ , \new_Sorter100|4270_ , \new_Sorter100|4271_ ,
    \new_Sorter100|4272_ , \new_Sorter100|4273_ , \new_Sorter100|4274_ ,
    \new_Sorter100|4275_ , \new_Sorter100|4276_ , \new_Sorter100|4277_ ,
    \new_Sorter100|4278_ , \new_Sorter100|4279_ , \new_Sorter100|4280_ ,
    \new_Sorter100|4281_ , \new_Sorter100|4282_ , \new_Sorter100|4283_ ,
    \new_Sorter100|4284_ , \new_Sorter100|4285_ , \new_Sorter100|4286_ ,
    \new_Sorter100|4287_ , \new_Sorter100|4288_ , \new_Sorter100|4289_ ,
    \new_Sorter100|4290_ , \new_Sorter100|4291_ , \new_Sorter100|4292_ ,
    \new_Sorter100|4293_ , \new_Sorter100|4294_ , \new_Sorter100|4295_ ,
    \new_Sorter100|4296_ , \new_Sorter100|4297_ , \new_Sorter100|4298_ ,
    \new_Sorter100|4299_ , \new_Sorter100|4300_ , \new_Sorter100|4399_ ,
    \new_Sorter100|4301_ , \new_Sorter100|4302_ , \new_Sorter100|4303_ ,
    \new_Sorter100|4304_ , \new_Sorter100|4305_ , \new_Sorter100|4306_ ,
    \new_Sorter100|4307_ , \new_Sorter100|4308_ , \new_Sorter100|4309_ ,
    \new_Sorter100|4310_ , \new_Sorter100|4311_ , \new_Sorter100|4312_ ,
    \new_Sorter100|4313_ , \new_Sorter100|4314_ , \new_Sorter100|4315_ ,
    \new_Sorter100|4316_ , \new_Sorter100|4317_ , \new_Sorter100|4318_ ,
    \new_Sorter100|4319_ , \new_Sorter100|4320_ , \new_Sorter100|4321_ ,
    \new_Sorter100|4322_ , \new_Sorter100|4323_ , \new_Sorter100|4324_ ,
    \new_Sorter100|4325_ , \new_Sorter100|4326_ , \new_Sorter100|4327_ ,
    \new_Sorter100|4328_ , \new_Sorter100|4329_ , \new_Sorter100|4330_ ,
    \new_Sorter100|4331_ , \new_Sorter100|4332_ , \new_Sorter100|4333_ ,
    \new_Sorter100|4334_ , \new_Sorter100|4335_ , \new_Sorter100|4336_ ,
    \new_Sorter100|4337_ , \new_Sorter100|4338_ , \new_Sorter100|4339_ ,
    \new_Sorter100|4340_ , \new_Sorter100|4341_ , \new_Sorter100|4342_ ,
    \new_Sorter100|4343_ , \new_Sorter100|4344_ , \new_Sorter100|4345_ ,
    \new_Sorter100|4346_ , \new_Sorter100|4347_ , \new_Sorter100|4348_ ,
    \new_Sorter100|4349_ , \new_Sorter100|4350_ , \new_Sorter100|4351_ ,
    \new_Sorter100|4352_ , \new_Sorter100|4353_ , \new_Sorter100|4354_ ,
    \new_Sorter100|4355_ , \new_Sorter100|4356_ , \new_Sorter100|4357_ ,
    \new_Sorter100|4358_ , \new_Sorter100|4359_ , \new_Sorter100|4360_ ,
    \new_Sorter100|4361_ , \new_Sorter100|4362_ , \new_Sorter100|4363_ ,
    \new_Sorter100|4364_ , \new_Sorter100|4365_ , \new_Sorter100|4366_ ,
    \new_Sorter100|4367_ , \new_Sorter100|4368_ , \new_Sorter100|4369_ ,
    \new_Sorter100|4370_ , \new_Sorter100|4371_ , \new_Sorter100|4372_ ,
    \new_Sorter100|4373_ , \new_Sorter100|4374_ , \new_Sorter100|4375_ ,
    \new_Sorter100|4376_ , \new_Sorter100|4377_ , \new_Sorter100|4378_ ,
    \new_Sorter100|4379_ , \new_Sorter100|4380_ , \new_Sorter100|4381_ ,
    \new_Sorter100|4382_ , \new_Sorter100|4383_ , \new_Sorter100|4384_ ,
    \new_Sorter100|4385_ , \new_Sorter100|4386_ , \new_Sorter100|4387_ ,
    \new_Sorter100|4388_ , \new_Sorter100|4389_ , \new_Sorter100|4390_ ,
    \new_Sorter100|4391_ , \new_Sorter100|4392_ , \new_Sorter100|4393_ ,
    \new_Sorter100|4394_ , \new_Sorter100|4395_ , \new_Sorter100|4396_ ,
    \new_Sorter100|4397_ , \new_Sorter100|4398_ , \new_Sorter100|4400_ ,
    \new_Sorter100|4401_ , \new_Sorter100|4402_ , \new_Sorter100|4403_ ,
    \new_Sorter100|4404_ , \new_Sorter100|4405_ , \new_Sorter100|4406_ ,
    \new_Sorter100|4407_ , \new_Sorter100|4408_ , \new_Sorter100|4409_ ,
    \new_Sorter100|4410_ , \new_Sorter100|4411_ , \new_Sorter100|4412_ ,
    \new_Sorter100|4413_ , \new_Sorter100|4414_ , \new_Sorter100|4415_ ,
    \new_Sorter100|4416_ , \new_Sorter100|4417_ , \new_Sorter100|4418_ ,
    \new_Sorter100|4419_ , \new_Sorter100|4420_ , \new_Sorter100|4421_ ,
    \new_Sorter100|4422_ , \new_Sorter100|4423_ , \new_Sorter100|4424_ ,
    \new_Sorter100|4425_ , \new_Sorter100|4426_ , \new_Sorter100|4427_ ,
    \new_Sorter100|4428_ , \new_Sorter100|4429_ , \new_Sorter100|4430_ ,
    \new_Sorter100|4431_ , \new_Sorter100|4432_ , \new_Sorter100|4433_ ,
    \new_Sorter100|4434_ , \new_Sorter100|4435_ , \new_Sorter100|4436_ ,
    \new_Sorter100|4437_ , \new_Sorter100|4438_ , \new_Sorter100|4439_ ,
    \new_Sorter100|4440_ , \new_Sorter100|4441_ , \new_Sorter100|4442_ ,
    \new_Sorter100|4443_ , \new_Sorter100|4444_ , \new_Sorter100|4445_ ,
    \new_Sorter100|4446_ , \new_Sorter100|4447_ , \new_Sorter100|4448_ ,
    \new_Sorter100|4449_ , \new_Sorter100|4450_ , \new_Sorter100|4451_ ,
    \new_Sorter100|4452_ , \new_Sorter100|4453_ , \new_Sorter100|4454_ ,
    \new_Sorter100|4455_ , \new_Sorter100|4456_ , \new_Sorter100|4457_ ,
    \new_Sorter100|4458_ , \new_Sorter100|4459_ , \new_Sorter100|4460_ ,
    \new_Sorter100|4461_ , \new_Sorter100|4462_ , \new_Sorter100|4463_ ,
    \new_Sorter100|4464_ , \new_Sorter100|4465_ , \new_Sorter100|4466_ ,
    \new_Sorter100|4467_ , \new_Sorter100|4468_ , \new_Sorter100|4469_ ,
    \new_Sorter100|4470_ , \new_Sorter100|4471_ , \new_Sorter100|4472_ ,
    \new_Sorter100|4473_ , \new_Sorter100|4474_ , \new_Sorter100|4475_ ,
    \new_Sorter100|4476_ , \new_Sorter100|4477_ , \new_Sorter100|4478_ ,
    \new_Sorter100|4479_ , \new_Sorter100|4480_ , \new_Sorter100|4481_ ,
    \new_Sorter100|4482_ , \new_Sorter100|4483_ , \new_Sorter100|4484_ ,
    \new_Sorter100|4485_ , \new_Sorter100|4486_ , \new_Sorter100|4487_ ,
    \new_Sorter100|4488_ , \new_Sorter100|4489_ , \new_Sorter100|4490_ ,
    \new_Sorter100|4491_ , \new_Sorter100|4492_ , \new_Sorter100|4493_ ,
    \new_Sorter100|4494_ , \new_Sorter100|4495_ , \new_Sorter100|4496_ ,
    \new_Sorter100|4497_ , \new_Sorter100|4498_ , \new_Sorter100|4499_ ,
    \new_Sorter100|4500_ , \new_Sorter100|4599_ , \new_Sorter100|4501_ ,
    \new_Sorter100|4502_ , \new_Sorter100|4503_ , \new_Sorter100|4504_ ,
    \new_Sorter100|4505_ , \new_Sorter100|4506_ , \new_Sorter100|4507_ ,
    \new_Sorter100|4508_ , \new_Sorter100|4509_ , \new_Sorter100|4510_ ,
    \new_Sorter100|4511_ , \new_Sorter100|4512_ , \new_Sorter100|4513_ ,
    \new_Sorter100|4514_ , \new_Sorter100|4515_ , \new_Sorter100|4516_ ,
    \new_Sorter100|4517_ , \new_Sorter100|4518_ , \new_Sorter100|4519_ ,
    \new_Sorter100|4520_ , \new_Sorter100|4521_ , \new_Sorter100|4522_ ,
    \new_Sorter100|4523_ , \new_Sorter100|4524_ , \new_Sorter100|4525_ ,
    \new_Sorter100|4526_ , \new_Sorter100|4527_ , \new_Sorter100|4528_ ,
    \new_Sorter100|4529_ , \new_Sorter100|4530_ , \new_Sorter100|4531_ ,
    \new_Sorter100|4532_ , \new_Sorter100|4533_ , \new_Sorter100|4534_ ,
    \new_Sorter100|4535_ , \new_Sorter100|4536_ , \new_Sorter100|4537_ ,
    \new_Sorter100|4538_ , \new_Sorter100|4539_ , \new_Sorter100|4540_ ,
    \new_Sorter100|4541_ , \new_Sorter100|4542_ , \new_Sorter100|4543_ ,
    \new_Sorter100|4544_ , \new_Sorter100|4545_ , \new_Sorter100|4546_ ,
    \new_Sorter100|4547_ , \new_Sorter100|4548_ , \new_Sorter100|4549_ ,
    \new_Sorter100|4550_ , \new_Sorter100|4551_ , \new_Sorter100|4552_ ,
    \new_Sorter100|4553_ , \new_Sorter100|4554_ , \new_Sorter100|4555_ ,
    \new_Sorter100|4556_ , \new_Sorter100|4557_ , \new_Sorter100|4558_ ,
    \new_Sorter100|4559_ , \new_Sorter100|4560_ , \new_Sorter100|4561_ ,
    \new_Sorter100|4562_ , \new_Sorter100|4563_ , \new_Sorter100|4564_ ,
    \new_Sorter100|4565_ , \new_Sorter100|4566_ , \new_Sorter100|4567_ ,
    \new_Sorter100|4568_ , \new_Sorter100|4569_ , \new_Sorter100|4570_ ,
    \new_Sorter100|4571_ , \new_Sorter100|4572_ , \new_Sorter100|4573_ ,
    \new_Sorter100|4574_ , \new_Sorter100|4575_ , \new_Sorter100|4576_ ,
    \new_Sorter100|4577_ , \new_Sorter100|4578_ , \new_Sorter100|4579_ ,
    \new_Sorter100|4580_ , \new_Sorter100|4581_ , \new_Sorter100|4582_ ,
    \new_Sorter100|4583_ , \new_Sorter100|4584_ , \new_Sorter100|4585_ ,
    \new_Sorter100|4586_ , \new_Sorter100|4587_ , \new_Sorter100|4588_ ,
    \new_Sorter100|4589_ , \new_Sorter100|4590_ , \new_Sorter100|4591_ ,
    \new_Sorter100|4592_ , \new_Sorter100|4593_ , \new_Sorter100|4594_ ,
    \new_Sorter100|4595_ , \new_Sorter100|4596_ , \new_Sorter100|4597_ ,
    \new_Sorter100|4598_ , \new_Sorter100|4600_ , \new_Sorter100|4601_ ,
    \new_Sorter100|4602_ , \new_Sorter100|4603_ , \new_Sorter100|4604_ ,
    \new_Sorter100|4605_ , \new_Sorter100|4606_ , \new_Sorter100|4607_ ,
    \new_Sorter100|4608_ , \new_Sorter100|4609_ , \new_Sorter100|4610_ ,
    \new_Sorter100|4611_ , \new_Sorter100|4612_ , \new_Sorter100|4613_ ,
    \new_Sorter100|4614_ , \new_Sorter100|4615_ , \new_Sorter100|4616_ ,
    \new_Sorter100|4617_ , \new_Sorter100|4618_ , \new_Sorter100|4619_ ,
    \new_Sorter100|4620_ , \new_Sorter100|4621_ , \new_Sorter100|4622_ ,
    \new_Sorter100|4623_ , \new_Sorter100|4624_ , \new_Sorter100|4625_ ,
    \new_Sorter100|4626_ , \new_Sorter100|4627_ , \new_Sorter100|4628_ ,
    \new_Sorter100|4629_ , \new_Sorter100|4630_ , \new_Sorter100|4631_ ,
    \new_Sorter100|4632_ , \new_Sorter100|4633_ , \new_Sorter100|4634_ ,
    \new_Sorter100|4635_ , \new_Sorter100|4636_ , \new_Sorter100|4637_ ,
    \new_Sorter100|4638_ , \new_Sorter100|4639_ , \new_Sorter100|4640_ ,
    \new_Sorter100|4641_ , \new_Sorter100|4642_ , \new_Sorter100|4643_ ,
    \new_Sorter100|4644_ , \new_Sorter100|4645_ , \new_Sorter100|4646_ ,
    \new_Sorter100|4647_ , \new_Sorter100|4648_ , \new_Sorter100|4649_ ,
    \new_Sorter100|4650_ , \new_Sorter100|4651_ , \new_Sorter100|4652_ ,
    \new_Sorter100|4653_ , \new_Sorter100|4654_ , \new_Sorter100|4655_ ,
    \new_Sorter100|4656_ , \new_Sorter100|4657_ , \new_Sorter100|4658_ ,
    \new_Sorter100|4659_ , \new_Sorter100|4660_ , \new_Sorter100|4661_ ,
    \new_Sorter100|4662_ , \new_Sorter100|4663_ , \new_Sorter100|4664_ ,
    \new_Sorter100|4665_ , \new_Sorter100|4666_ , \new_Sorter100|4667_ ,
    \new_Sorter100|4668_ , \new_Sorter100|4669_ , \new_Sorter100|4670_ ,
    \new_Sorter100|4671_ , \new_Sorter100|4672_ , \new_Sorter100|4673_ ,
    \new_Sorter100|4674_ , \new_Sorter100|4675_ , \new_Sorter100|4676_ ,
    \new_Sorter100|4677_ , \new_Sorter100|4678_ , \new_Sorter100|4679_ ,
    \new_Sorter100|4680_ , \new_Sorter100|4681_ , \new_Sorter100|4682_ ,
    \new_Sorter100|4683_ , \new_Sorter100|4684_ , \new_Sorter100|4685_ ,
    \new_Sorter100|4686_ , \new_Sorter100|4687_ , \new_Sorter100|4688_ ,
    \new_Sorter100|4689_ , \new_Sorter100|4690_ , \new_Sorter100|4691_ ,
    \new_Sorter100|4692_ , \new_Sorter100|4693_ , \new_Sorter100|4694_ ,
    \new_Sorter100|4695_ , \new_Sorter100|4696_ , \new_Sorter100|4697_ ,
    \new_Sorter100|4698_ , \new_Sorter100|4699_ , \new_Sorter100|4700_ ,
    \new_Sorter100|4799_ , \new_Sorter100|4701_ , \new_Sorter100|4702_ ,
    \new_Sorter100|4703_ , \new_Sorter100|4704_ , \new_Sorter100|4705_ ,
    \new_Sorter100|4706_ , \new_Sorter100|4707_ , \new_Sorter100|4708_ ,
    \new_Sorter100|4709_ , \new_Sorter100|4710_ , \new_Sorter100|4711_ ,
    \new_Sorter100|4712_ , \new_Sorter100|4713_ , \new_Sorter100|4714_ ,
    \new_Sorter100|4715_ , \new_Sorter100|4716_ , \new_Sorter100|4717_ ,
    \new_Sorter100|4718_ , \new_Sorter100|4719_ , \new_Sorter100|4720_ ,
    \new_Sorter100|4721_ , \new_Sorter100|4722_ , \new_Sorter100|4723_ ,
    \new_Sorter100|4724_ , \new_Sorter100|4725_ , \new_Sorter100|4726_ ,
    \new_Sorter100|4727_ , \new_Sorter100|4728_ , \new_Sorter100|4729_ ,
    \new_Sorter100|4730_ , \new_Sorter100|4731_ , \new_Sorter100|4732_ ,
    \new_Sorter100|4733_ , \new_Sorter100|4734_ , \new_Sorter100|4735_ ,
    \new_Sorter100|4736_ , \new_Sorter100|4737_ , \new_Sorter100|4738_ ,
    \new_Sorter100|4739_ , \new_Sorter100|4740_ , \new_Sorter100|4741_ ,
    \new_Sorter100|4742_ , \new_Sorter100|4743_ , \new_Sorter100|4744_ ,
    \new_Sorter100|4745_ , \new_Sorter100|4746_ , \new_Sorter100|4747_ ,
    \new_Sorter100|4748_ , \new_Sorter100|4749_ , \new_Sorter100|4750_ ,
    \new_Sorter100|4751_ , \new_Sorter100|4752_ , \new_Sorter100|4753_ ,
    \new_Sorter100|4754_ , \new_Sorter100|4755_ , \new_Sorter100|4756_ ,
    \new_Sorter100|4757_ , \new_Sorter100|4758_ , \new_Sorter100|4759_ ,
    \new_Sorter100|4760_ , \new_Sorter100|4761_ , \new_Sorter100|4762_ ,
    \new_Sorter100|4763_ , \new_Sorter100|4764_ , \new_Sorter100|4765_ ,
    \new_Sorter100|4766_ , \new_Sorter100|4767_ , \new_Sorter100|4768_ ,
    \new_Sorter100|4769_ , \new_Sorter100|4770_ , \new_Sorter100|4771_ ,
    \new_Sorter100|4772_ , \new_Sorter100|4773_ , \new_Sorter100|4774_ ,
    \new_Sorter100|4775_ , \new_Sorter100|4776_ , \new_Sorter100|4777_ ,
    \new_Sorter100|4778_ , \new_Sorter100|4779_ , \new_Sorter100|4780_ ,
    \new_Sorter100|4781_ , \new_Sorter100|4782_ , \new_Sorter100|4783_ ,
    \new_Sorter100|4784_ , \new_Sorter100|4785_ , \new_Sorter100|4786_ ,
    \new_Sorter100|4787_ , \new_Sorter100|4788_ , \new_Sorter100|4789_ ,
    \new_Sorter100|4790_ , \new_Sorter100|4791_ , \new_Sorter100|4792_ ,
    \new_Sorter100|4793_ , \new_Sorter100|4794_ , \new_Sorter100|4795_ ,
    \new_Sorter100|4796_ , \new_Sorter100|4797_ , \new_Sorter100|4798_ ,
    \new_Sorter100|4800_ , \new_Sorter100|4801_ , \new_Sorter100|4802_ ,
    \new_Sorter100|4803_ , \new_Sorter100|4804_ , \new_Sorter100|4805_ ,
    \new_Sorter100|4806_ , \new_Sorter100|4807_ , \new_Sorter100|4808_ ,
    \new_Sorter100|4809_ , \new_Sorter100|4810_ , \new_Sorter100|4811_ ,
    \new_Sorter100|4812_ , \new_Sorter100|4813_ , \new_Sorter100|4814_ ,
    \new_Sorter100|4815_ , \new_Sorter100|4816_ , \new_Sorter100|4817_ ,
    \new_Sorter100|4818_ , \new_Sorter100|4819_ , \new_Sorter100|4820_ ,
    \new_Sorter100|4821_ , \new_Sorter100|4822_ , \new_Sorter100|4823_ ,
    \new_Sorter100|4824_ , \new_Sorter100|4825_ , \new_Sorter100|4826_ ,
    \new_Sorter100|4827_ , \new_Sorter100|4828_ , \new_Sorter100|4829_ ,
    \new_Sorter100|4830_ , \new_Sorter100|4831_ , \new_Sorter100|4832_ ,
    \new_Sorter100|4833_ , \new_Sorter100|4834_ , \new_Sorter100|4835_ ,
    \new_Sorter100|4836_ , \new_Sorter100|4837_ , \new_Sorter100|4838_ ,
    \new_Sorter100|4839_ , \new_Sorter100|4840_ , \new_Sorter100|4841_ ,
    \new_Sorter100|4842_ , \new_Sorter100|4843_ , \new_Sorter100|4844_ ,
    \new_Sorter100|4845_ , \new_Sorter100|4846_ , \new_Sorter100|4847_ ,
    \new_Sorter100|4848_ , \new_Sorter100|4849_ , \new_Sorter100|4850_ ,
    \new_Sorter100|4851_ , \new_Sorter100|4852_ , \new_Sorter100|4853_ ,
    \new_Sorter100|4854_ , \new_Sorter100|4855_ , \new_Sorter100|4856_ ,
    \new_Sorter100|4857_ , \new_Sorter100|4858_ , \new_Sorter100|4859_ ,
    \new_Sorter100|4860_ , \new_Sorter100|4861_ , \new_Sorter100|4862_ ,
    \new_Sorter100|4863_ , \new_Sorter100|4864_ , \new_Sorter100|4865_ ,
    \new_Sorter100|4866_ , \new_Sorter100|4867_ , \new_Sorter100|4868_ ,
    \new_Sorter100|4869_ , \new_Sorter100|4870_ , \new_Sorter100|4871_ ,
    \new_Sorter100|4872_ , \new_Sorter100|4873_ , \new_Sorter100|4874_ ,
    \new_Sorter100|4875_ , \new_Sorter100|4876_ , \new_Sorter100|4877_ ,
    \new_Sorter100|4878_ , \new_Sorter100|4879_ , \new_Sorter100|4880_ ,
    \new_Sorter100|4881_ , \new_Sorter100|4882_ , \new_Sorter100|4883_ ,
    \new_Sorter100|4884_ , \new_Sorter100|4885_ , \new_Sorter100|4886_ ,
    \new_Sorter100|4887_ , \new_Sorter100|4888_ , \new_Sorter100|4889_ ,
    \new_Sorter100|4890_ , \new_Sorter100|4891_ , \new_Sorter100|4892_ ,
    \new_Sorter100|4893_ , \new_Sorter100|4894_ , \new_Sorter100|4895_ ,
    \new_Sorter100|4896_ , \new_Sorter100|4897_ , \new_Sorter100|4898_ ,
    \new_Sorter100|4899_ , \new_Sorter100|4900_ , \new_Sorter100|4999_ ,
    \new_Sorter100|4901_ , \new_Sorter100|4902_ , \new_Sorter100|4903_ ,
    \new_Sorter100|4904_ , \new_Sorter100|4905_ , \new_Sorter100|4906_ ,
    \new_Sorter100|4907_ , \new_Sorter100|4908_ , \new_Sorter100|4909_ ,
    \new_Sorter100|4910_ , \new_Sorter100|4911_ , \new_Sorter100|4912_ ,
    \new_Sorter100|4913_ , \new_Sorter100|4914_ , \new_Sorter100|4915_ ,
    \new_Sorter100|4916_ , \new_Sorter100|4917_ , \new_Sorter100|4918_ ,
    \new_Sorter100|4919_ , \new_Sorter100|4920_ , \new_Sorter100|4921_ ,
    \new_Sorter100|4922_ , \new_Sorter100|4923_ , \new_Sorter100|4924_ ,
    \new_Sorter100|4925_ , \new_Sorter100|4926_ , \new_Sorter100|4927_ ,
    \new_Sorter100|4928_ , \new_Sorter100|4929_ , \new_Sorter100|4930_ ,
    \new_Sorter100|4931_ , \new_Sorter100|4932_ , \new_Sorter100|4933_ ,
    \new_Sorter100|4934_ , \new_Sorter100|4935_ , \new_Sorter100|4936_ ,
    \new_Sorter100|4937_ , \new_Sorter100|4938_ , \new_Sorter100|4939_ ,
    \new_Sorter100|4940_ , \new_Sorter100|4941_ , \new_Sorter100|4942_ ,
    \new_Sorter100|4943_ , \new_Sorter100|4944_ , \new_Sorter100|4945_ ,
    \new_Sorter100|4946_ , \new_Sorter100|4947_ , \new_Sorter100|4948_ ,
    \new_Sorter100|4949_ , \new_Sorter100|4950_ , \new_Sorter100|4951_ ,
    \new_Sorter100|4952_ , \new_Sorter100|4953_ , \new_Sorter100|4954_ ,
    \new_Sorter100|4955_ , \new_Sorter100|4956_ , \new_Sorter100|4957_ ,
    \new_Sorter100|4958_ , \new_Sorter100|4959_ , \new_Sorter100|4960_ ,
    \new_Sorter100|4961_ , \new_Sorter100|4962_ , \new_Sorter100|4963_ ,
    \new_Sorter100|4964_ , \new_Sorter100|4965_ , \new_Sorter100|4966_ ,
    \new_Sorter100|4967_ , \new_Sorter100|4968_ , \new_Sorter100|4969_ ,
    \new_Sorter100|4970_ , \new_Sorter100|4971_ , \new_Sorter100|4972_ ,
    \new_Sorter100|4973_ , \new_Sorter100|4974_ , \new_Sorter100|4975_ ,
    \new_Sorter100|4976_ , \new_Sorter100|4977_ , \new_Sorter100|4978_ ,
    \new_Sorter100|4979_ , \new_Sorter100|4980_ , \new_Sorter100|4981_ ,
    \new_Sorter100|4982_ , \new_Sorter100|4983_ , \new_Sorter100|4984_ ,
    \new_Sorter100|4985_ , \new_Sorter100|4986_ , \new_Sorter100|4987_ ,
    \new_Sorter100|4988_ , \new_Sorter100|4989_ , \new_Sorter100|4990_ ,
    \new_Sorter100|4991_ , \new_Sorter100|4992_ , \new_Sorter100|4993_ ,
    \new_Sorter100|4994_ , \new_Sorter100|4995_ , \new_Sorter100|4996_ ,
    \new_Sorter100|4997_ , \new_Sorter100|4998_ , \new_Sorter100|5000_ ,
    \new_Sorter100|5001_ , \new_Sorter100|5002_ , \new_Sorter100|5003_ ,
    \new_Sorter100|5004_ , \new_Sorter100|5005_ , \new_Sorter100|5006_ ,
    \new_Sorter100|5007_ , \new_Sorter100|5008_ , \new_Sorter100|5009_ ,
    \new_Sorter100|5010_ , \new_Sorter100|5011_ , \new_Sorter100|5012_ ,
    \new_Sorter100|5013_ , \new_Sorter100|5014_ , \new_Sorter100|5015_ ,
    \new_Sorter100|5016_ , \new_Sorter100|5017_ , \new_Sorter100|5018_ ,
    \new_Sorter100|5019_ , \new_Sorter100|5020_ , \new_Sorter100|5021_ ,
    \new_Sorter100|5022_ , \new_Sorter100|5023_ , \new_Sorter100|5024_ ,
    \new_Sorter100|5025_ , \new_Sorter100|5026_ , \new_Sorter100|5027_ ,
    \new_Sorter100|5028_ , \new_Sorter100|5029_ , \new_Sorter100|5030_ ,
    \new_Sorter100|5031_ , \new_Sorter100|5032_ , \new_Sorter100|5033_ ,
    \new_Sorter100|5034_ , \new_Sorter100|5035_ , \new_Sorter100|5036_ ,
    \new_Sorter100|5037_ , \new_Sorter100|5038_ , \new_Sorter100|5039_ ,
    \new_Sorter100|5040_ , \new_Sorter100|5041_ , \new_Sorter100|5042_ ,
    \new_Sorter100|5043_ , \new_Sorter100|5044_ , \new_Sorter100|5045_ ,
    \new_Sorter100|5046_ , \new_Sorter100|5047_ , \new_Sorter100|5048_ ,
    \new_Sorter100|5049_ , \new_Sorter100|5050_ , \new_Sorter100|5051_ ,
    \new_Sorter100|5052_ , \new_Sorter100|5053_ , \new_Sorter100|5054_ ,
    \new_Sorter100|5055_ , \new_Sorter100|5056_ , \new_Sorter100|5057_ ,
    \new_Sorter100|5058_ , \new_Sorter100|5059_ , \new_Sorter100|5060_ ,
    \new_Sorter100|5061_ , \new_Sorter100|5062_ , \new_Sorter100|5063_ ,
    \new_Sorter100|5064_ , \new_Sorter100|5065_ , \new_Sorter100|5066_ ,
    \new_Sorter100|5067_ , \new_Sorter100|5068_ , \new_Sorter100|5069_ ,
    \new_Sorter100|5070_ , \new_Sorter100|5071_ , \new_Sorter100|5072_ ,
    \new_Sorter100|5073_ , \new_Sorter100|5074_ , \new_Sorter100|5075_ ,
    \new_Sorter100|5076_ , \new_Sorter100|5077_ , \new_Sorter100|5078_ ,
    \new_Sorter100|5079_ , \new_Sorter100|5080_ , \new_Sorter100|5081_ ,
    \new_Sorter100|5082_ , \new_Sorter100|5083_ , \new_Sorter100|5084_ ,
    \new_Sorter100|5085_ , \new_Sorter100|5086_ , \new_Sorter100|5087_ ,
    \new_Sorter100|5088_ , \new_Sorter100|5089_ , \new_Sorter100|5090_ ,
    \new_Sorter100|5091_ , \new_Sorter100|5092_ , \new_Sorter100|5093_ ,
    \new_Sorter100|5094_ , \new_Sorter100|5095_ , \new_Sorter100|5096_ ,
    \new_Sorter100|5097_ , \new_Sorter100|5098_ , \new_Sorter100|5099_ ,
    \new_Sorter100|5100_ , \new_Sorter100|5199_ , \new_Sorter100|5101_ ,
    \new_Sorter100|5102_ , \new_Sorter100|5103_ , \new_Sorter100|5104_ ,
    \new_Sorter100|5105_ , \new_Sorter100|5106_ , \new_Sorter100|5107_ ,
    \new_Sorter100|5108_ , \new_Sorter100|5109_ , \new_Sorter100|5110_ ,
    \new_Sorter100|5111_ , \new_Sorter100|5112_ , \new_Sorter100|5113_ ,
    \new_Sorter100|5114_ , \new_Sorter100|5115_ , \new_Sorter100|5116_ ,
    \new_Sorter100|5117_ , \new_Sorter100|5118_ , \new_Sorter100|5119_ ,
    \new_Sorter100|5120_ , \new_Sorter100|5121_ , \new_Sorter100|5122_ ,
    \new_Sorter100|5123_ , \new_Sorter100|5124_ , \new_Sorter100|5125_ ,
    \new_Sorter100|5126_ , \new_Sorter100|5127_ , \new_Sorter100|5128_ ,
    \new_Sorter100|5129_ , \new_Sorter100|5130_ , \new_Sorter100|5131_ ,
    \new_Sorter100|5132_ , \new_Sorter100|5133_ , \new_Sorter100|5134_ ,
    \new_Sorter100|5135_ , \new_Sorter100|5136_ , \new_Sorter100|5137_ ,
    \new_Sorter100|5138_ , \new_Sorter100|5139_ , \new_Sorter100|5140_ ,
    \new_Sorter100|5141_ , \new_Sorter100|5142_ , \new_Sorter100|5143_ ,
    \new_Sorter100|5144_ , \new_Sorter100|5145_ , \new_Sorter100|5146_ ,
    \new_Sorter100|5147_ , \new_Sorter100|5148_ , \new_Sorter100|5149_ ,
    \new_Sorter100|5150_ , \new_Sorter100|5151_ , \new_Sorter100|5152_ ,
    \new_Sorter100|5153_ , \new_Sorter100|5154_ , \new_Sorter100|5155_ ,
    \new_Sorter100|5156_ , \new_Sorter100|5157_ , \new_Sorter100|5158_ ,
    \new_Sorter100|5159_ , \new_Sorter100|5160_ , \new_Sorter100|5161_ ,
    \new_Sorter100|5162_ , \new_Sorter100|5163_ , \new_Sorter100|5164_ ,
    \new_Sorter100|5165_ , \new_Sorter100|5166_ , \new_Sorter100|5167_ ,
    \new_Sorter100|5168_ , \new_Sorter100|5169_ , \new_Sorter100|5170_ ,
    \new_Sorter100|5171_ , \new_Sorter100|5172_ , \new_Sorter100|5173_ ,
    \new_Sorter100|5174_ , \new_Sorter100|5175_ , \new_Sorter100|5176_ ,
    \new_Sorter100|5177_ , \new_Sorter100|5178_ , \new_Sorter100|5179_ ,
    \new_Sorter100|5180_ , \new_Sorter100|5181_ , \new_Sorter100|5182_ ,
    \new_Sorter100|5183_ , \new_Sorter100|5184_ , \new_Sorter100|5185_ ,
    \new_Sorter100|5186_ , \new_Sorter100|5187_ , \new_Sorter100|5188_ ,
    \new_Sorter100|5189_ , \new_Sorter100|5190_ , \new_Sorter100|5191_ ,
    \new_Sorter100|5192_ , \new_Sorter100|5193_ , \new_Sorter100|5194_ ,
    \new_Sorter100|5195_ , \new_Sorter100|5196_ , \new_Sorter100|5197_ ,
    \new_Sorter100|5198_ , \new_Sorter100|5200_ , \new_Sorter100|5201_ ,
    \new_Sorter100|5202_ , \new_Sorter100|5203_ , \new_Sorter100|5204_ ,
    \new_Sorter100|5205_ , \new_Sorter100|5206_ , \new_Sorter100|5207_ ,
    \new_Sorter100|5208_ , \new_Sorter100|5209_ , \new_Sorter100|5210_ ,
    \new_Sorter100|5211_ , \new_Sorter100|5212_ , \new_Sorter100|5213_ ,
    \new_Sorter100|5214_ , \new_Sorter100|5215_ , \new_Sorter100|5216_ ,
    \new_Sorter100|5217_ , \new_Sorter100|5218_ , \new_Sorter100|5219_ ,
    \new_Sorter100|5220_ , \new_Sorter100|5221_ , \new_Sorter100|5222_ ,
    \new_Sorter100|5223_ , \new_Sorter100|5224_ , \new_Sorter100|5225_ ,
    \new_Sorter100|5226_ , \new_Sorter100|5227_ , \new_Sorter100|5228_ ,
    \new_Sorter100|5229_ , \new_Sorter100|5230_ , \new_Sorter100|5231_ ,
    \new_Sorter100|5232_ , \new_Sorter100|5233_ , \new_Sorter100|5234_ ,
    \new_Sorter100|5235_ , \new_Sorter100|5236_ , \new_Sorter100|5237_ ,
    \new_Sorter100|5238_ , \new_Sorter100|5239_ , \new_Sorter100|5240_ ,
    \new_Sorter100|5241_ , \new_Sorter100|5242_ , \new_Sorter100|5243_ ,
    \new_Sorter100|5244_ , \new_Sorter100|5245_ , \new_Sorter100|5246_ ,
    \new_Sorter100|5247_ , \new_Sorter100|5248_ , \new_Sorter100|5249_ ,
    \new_Sorter100|5250_ , \new_Sorter100|5251_ , \new_Sorter100|5252_ ,
    \new_Sorter100|5253_ , \new_Sorter100|5254_ , \new_Sorter100|5255_ ,
    \new_Sorter100|5256_ , \new_Sorter100|5257_ , \new_Sorter100|5258_ ,
    \new_Sorter100|5259_ , \new_Sorter100|5260_ , \new_Sorter100|5261_ ,
    \new_Sorter100|5262_ , \new_Sorter100|5263_ , \new_Sorter100|5264_ ,
    \new_Sorter100|5265_ , \new_Sorter100|5266_ , \new_Sorter100|5267_ ,
    \new_Sorter100|5268_ , \new_Sorter100|5269_ , \new_Sorter100|5270_ ,
    \new_Sorter100|5271_ , \new_Sorter100|5272_ , \new_Sorter100|5273_ ,
    \new_Sorter100|5274_ , \new_Sorter100|5275_ , \new_Sorter100|5276_ ,
    \new_Sorter100|5277_ , \new_Sorter100|5278_ , \new_Sorter100|5279_ ,
    \new_Sorter100|5280_ , \new_Sorter100|5281_ , \new_Sorter100|5282_ ,
    \new_Sorter100|5283_ , \new_Sorter100|5284_ , \new_Sorter100|5285_ ,
    \new_Sorter100|5286_ , \new_Sorter100|5287_ , \new_Sorter100|5288_ ,
    \new_Sorter100|5289_ , \new_Sorter100|5290_ , \new_Sorter100|5291_ ,
    \new_Sorter100|5292_ , \new_Sorter100|5293_ , \new_Sorter100|5294_ ,
    \new_Sorter100|5295_ , \new_Sorter100|5296_ , \new_Sorter100|5297_ ,
    \new_Sorter100|5298_ , \new_Sorter100|5299_ , \new_Sorter100|5300_ ,
    \new_Sorter100|5399_ , \new_Sorter100|5301_ , \new_Sorter100|5302_ ,
    \new_Sorter100|5303_ , \new_Sorter100|5304_ , \new_Sorter100|5305_ ,
    \new_Sorter100|5306_ , \new_Sorter100|5307_ , \new_Sorter100|5308_ ,
    \new_Sorter100|5309_ , \new_Sorter100|5310_ , \new_Sorter100|5311_ ,
    \new_Sorter100|5312_ , \new_Sorter100|5313_ , \new_Sorter100|5314_ ,
    \new_Sorter100|5315_ , \new_Sorter100|5316_ , \new_Sorter100|5317_ ,
    \new_Sorter100|5318_ , \new_Sorter100|5319_ , \new_Sorter100|5320_ ,
    \new_Sorter100|5321_ , \new_Sorter100|5322_ , \new_Sorter100|5323_ ,
    \new_Sorter100|5324_ , \new_Sorter100|5325_ , \new_Sorter100|5326_ ,
    \new_Sorter100|5327_ , \new_Sorter100|5328_ , \new_Sorter100|5329_ ,
    \new_Sorter100|5330_ , \new_Sorter100|5331_ , \new_Sorter100|5332_ ,
    \new_Sorter100|5333_ , \new_Sorter100|5334_ , \new_Sorter100|5335_ ,
    \new_Sorter100|5336_ , \new_Sorter100|5337_ , \new_Sorter100|5338_ ,
    \new_Sorter100|5339_ , \new_Sorter100|5340_ , \new_Sorter100|5341_ ,
    \new_Sorter100|5342_ , \new_Sorter100|5343_ , \new_Sorter100|5344_ ,
    \new_Sorter100|5345_ , \new_Sorter100|5346_ , \new_Sorter100|5347_ ,
    \new_Sorter100|5348_ , \new_Sorter100|5349_ , \new_Sorter100|5350_ ,
    \new_Sorter100|5351_ , \new_Sorter100|5352_ , \new_Sorter100|5353_ ,
    \new_Sorter100|5354_ , \new_Sorter100|5355_ , \new_Sorter100|5356_ ,
    \new_Sorter100|5357_ , \new_Sorter100|5358_ , \new_Sorter100|5359_ ,
    \new_Sorter100|5360_ , \new_Sorter100|5361_ , \new_Sorter100|5362_ ,
    \new_Sorter100|5363_ , \new_Sorter100|5364_ , \new_Sorter100|5365_ ,
    \new_Sorter100|5366_ , \new_Sorter100|5367_ , \new_Sorter100|5368_ ,
    \new_Sorter100|5369_ , \new_Sorter100|5370_ , \new_Sorter100|5371_ ,
    \new_Sorter100|5372_ , \new_Sorter100|5373_ , \new_Sorter100|5374_ ,
    \new_Sorter100|5375_ , \new_Sorter100|5376_ , \new_Sorter100|5377_ ,
    \new_Sorter100|5378_ , \new_Sorter100|5379_ , \new_Sorter100|5380_ ,
    \new_Sorter100|5381_ , \new_Sorter100|5382_ , \new_Sorter100|5383_ ,
    \new_Sorter100|5384_ , \new_Sorter100|5385_ , \new_Sorter100|5386_ ,
    \new_Sorter100|5387_ , \new_Sorter100|5388_ , \new_Sorter100|5389_ ,
    \new_Sorter100|5390_ , \new_Sorter100|5391_ , \new_Sorter100|5392_ ,
    \new_Sorter100|5393_ , \new_Sorter100|5394_ , \new_Sorter100|5395_ ,
    \new_Sorter100|5396_ , \new_Sorter100|5397_ , \new_Sorter100|5398_ ,
    \new_Sorter100|5400_ , \new_Sorter100|5401_ , \new_Sorter100|5402_ ,
    \new_Sorter100|5403_ , \new_Sorter100|5404_ , \new_Sorter100|5405_ ,
    \new_Sorter100|5406_ , \new_Sorter100|5407_ , \new_Sorter100|5408_ ,
    \new_Sorter100|5409_ , \new_Sorter100|5410_ , \new_Sorter100|5411_ ,
    \new_Sorter100|5412_ , \new_Sorter100|5413_ , \new_Sorter100|5414_ ,
    \new_Sorter100|5415_ , \new_Sorter100|5416_ , \new_Sorter100|5417_ ,
    \new_Sorter100|5418_ , \new_Sorter100|5419_ , \new_Sorter100|5420_ ,
    \new_Sorter100|5421_ , \new_Sorter100|5422_ , \new_Sorter100|5423_ ,
    \new_Sorter100|5424_ , \new_Sorter100|5425_ , \new_Sorter100|5426_ ,
    \new_Sorter100|5427_ , \new_Sorter100|5428_ , \new_Sorter100|5429_ ,
    \new_Sorter100|5430_ , \new_Sorter100|5431_ , \new_Sorter100|5432_ ,
    \new_Sorter100|5433_ , \new_Sorter100|5434_ , \new_Sorter100|5435_ ,
    \new_Sorter100|5436_ , \new_Sorter100|5437_ , \new_Sorter100|5438_ ,
    \new_Sorter100|5439_ , \new_Sorter100|5440_ , \new_Sorter100|5441_ ,
    \new_Sorter100|5442_ , \new_Sorter100|5443_ , \new_Sorter100|5444_ ,
    \new_Sorter100|5445_ , \new_Sorter100|5446_ , \new_Sorter100|5447_ ,
    \new_Sorter100|5448_ , \new_Sorter100|5449_ , \new_Sorter100|5450_ ,
    \new_Sorter100|5451_ , \new_Sorter100|5452_ , \new_Sorter100|5453_ ,
    \new_Sorter100|5454_ , \new_Sorter100|5455_ , \new_Sorter100|5456_ ,
    \new_Sorter100|5457_ , \new_Sorter100|5458_ , \new_Sorter100|5459_ ,
    \new_Sorter100|5460_ , \new_Sorter100|5461_ , \new_Sorter100|5462_ ,
    \new_Sorter100|5463_ , \new_Sorter100|5464_ , \new_Sorter100|5465_ ,
    \new_Sorter100|5466_ , \new_Sorter100|5467_ , \new_Sorter100|5468_ ,
    \new_Sorter100|5469_ , \new_Sorter100|5470_ , \new_Sorter100|5471_ ,
    \new_Sorter100|5472_ , \new_Sorter100|5473_ , \new_Sorter100|5474_ ,
    \new_Sorter100|5475_ , \new_Sorter100|5476_ , \new_Sorter100|5477_ ,
    \new_Sorter100|5478_ , \new_Sorter100|5479_ , \new_Sorter100|5480_ ,
    \new_Sorter100|5481_ , \new_Sorter100|5482_ , \new_Sorter100|5483_ ,
    \new_Sorter100|5484_ , \new_Sorter100|5485_ , \new_Sorter100|5486_ ,
    \new_Sorter100|5487_ , \new_Sorter100|5488_ , \new_Sorter100|5489_ ,
    \new_Sorter100|5490_ , \new_Sorter100|5491_ , \new_Sorter100|5492_ ,
    \new_Sorter100|5493_ , \new_Sorter100|5494_ , \new_Sorter100|5495_ ,
    \new_Sorter100|5496_ , \new_Sorter100|5497_ , \new_Sorter100|5498_ ,
    \new_Sorter100|5499_ , \new_Sorter100|5500_ , \new_Sorter100|5599_ ,
    \new_Sorter100|5501_ , \new_Sorter100|5502_ , \new_Sorter100|5503_ ,
    \new_Sorter100|5504_ , \new_Sorter100|5505_ , \new_Sorter100|5506_ ,
    \new_Sorter100|5507_ , \new_Sorter100|5508_ , \new_Sorter100|5509_ ,
    \new_Sorter100|5510_ , \new_Sorter100|5511_ , \new_Sorter100|5512_ ,
    \new_Sorter100|5513_ , \new_Sorter100|5514_ , \new_Sorter100|5515_ ,
    \new_Sorter100|5516_ , \new_Sorter100|5517_ , \new_Sorter100|5518_ ,
    \new_Sorter100|5519_ , \new_Sorter100|5520_ , \new_Sorter100|5521_ ,
    \new_Sorter100|5522_ , \new_Sorter100|5523_ , \new_Sorter100|5524_ ,
    \new_Sorter100|5525_ , \new_Sorter100|5526_ , \new_Sorter100|5527_ ,
    \new_Sorter100|5528_ , \new_Sorter100|5529_ , \new_Sorter100|5530_ ,
    \new_Sorter100|5531_ , \new_Sorter100|5532_ , \new_Sorter100|5533_ ,
    \new_Sorter100|5534_ , \new_Sorter100|5535_ , \new_Sorter100|5536_ ,
    \new_Sorter100|5537_ , \new_Sorter100|5538_ , \new_Sorter100|5539_ ,
    \new_Sorter100|5540_ , \new_Sorter100|5541_ , \new_Sorter100|5542_ ,
    \new_Sorter100|5543_ , \new_Sorter100|5544_ , \new_Sorter100|5545_ ,
    \new_Sorter100|5546_ , \new_Sorter100|5547_ , \new_Sorter100|5548_ ,
    \new_Sorter100|5549_ , \new_Sorter100|5550_ , \new_Sorter100|5551_ ,
    \new_Sorter100|5552_ , \new_Sorter100|5553_ , \new_Sorter100|5554_ ,
    \new_Sorter100|5555_ , \new_Sorter100|5556_ , \new_Sorter100|5557_ ,
    \new_Sorter100|5558_ , \new_Sorter100|5559_ , \new_Sorter100|5560_ ,
    \new_Sorter100|5561_ , \new_Sorter100|5562_ , \new_Sorter100|5563_ ,
    \new_Sorter100|5564_ , \new_Sorter100|5565_ , \new_Sorter100|5566_ ,
    \new_Sorter100|5567_ , \new_Sorter100|5568_ , \new_Sorter100|5569_ ,
    \new_Sorter100|5570_ , \new_Sorter100|5571_ , \new_Sorter100|5572_ ,
    \new_Sorter100|5573_ , \new_Sorter100|5574_ , \new_Sorter100|5575_ ,
    \new_Sorter100|5576_ , \new_Sorter100|5577_ , \new_Sorter100|5578_ ,
    \new_Sorter100|5579_ , \new_Sorter100|5580_ , \new_Sorter100|5581_ ,
    \new_Sorter100|5582_ , \new_Sorter100|5583_ , \new_Sorter100|5584_ ,
    \new_Sorter100|5585_ , \new_Sorter100|5586_ , \new_Sorter100|5587_ ,
    \new_Sorter100|5588_ , \new_Sorter100|5589_ , \new_Sorter100|5590_ ,
    \new_Sorter100|5591_ , \new_Sorter100|5592_ , \new_Sorter100|5593_ ,
    \new_Sorter100|5594_ , \new_Sorter100|5595_ , \new_Sorter100|5596_ ,
    \new_Sorter100|5597_ , \new_Sorter100|5598_ , \new_Sorter100|5600_ ,
    \new_Sorter100|5601_ , \new_Sorter100|5602_ , \new_Sorter100|5603_ ,
    \new_Sorter100|5604_ , \new_Sorter100|5605_ , \new_Sorter100|5606_ ,
    \new_Sorter100|5607_ , \new_Sorter100|5608_ , \new_Sorter100|5609_ ,
    \new_Sorter100|5610_ , \new_Sorter100|5611_ , \new_Sorter100|5612_ ,
    \new_Sorter100|5613_ , \new_Sorter100|5614_ , \new_Sorter100|5615_ ,
    \new_Sorter100|5616_ , \new_Sorter100|5617_ , \new_Sorter100|5618_ ,
    \new_Sorter100|5619_ , \new_Sorter100|5620_ , \new_Sorter100|5621_ ,
    \new_Sorter100|5622_ , \new_Sorter100|5623_ , \new_Sorter100|5624_ ,
    \new_Sorter100|5625_ , \new_Sorter100|5626_ , \new_Sorter100|5627_ ,
    \new_Sorter100|5628_ , \new_Sorter100|5629_ , \new_Sorter100|5630_ ,
    \new_Sorter100|5631_ , \new_Sorter100|5632_ , \new_Sorter100|5633_ ,
    \new_Sorter100|5634_ , \new_Sorter100|5635_ , \new_Sorter100|5636_ ,
    \new_Sorter100|5637_ , \new_Sorter100|5638_ , \new_Sorter100|5639_ ,
    \new_Sorter100|5640_ , \new_Sorter100|5641_ , \new_Sorter100|5642_ ,
    \new_Sorter100|5643_ , \new_Sorter100|5644_ , \new_Sorter100|5645_ ,
    \new_Sorter100|5646_ , \new_Sorter100|5647_ , \new_Sorter100|5648_ ,
    \new_Sorter100|5649_ , \new_Sorter100|5650_ , \new_Sorter100|5651_ ,
    \new_Sorter100|5652_ , \new_Sorter100|5653_ , \new_Sorter100|5654_ ,
    \new_Sorter100|5655_ , \new_Sorter100|5656_ , \new_Sorter100|5657_ ,
    \new_Sorter100|5658_ , \new_Sorter100|5659_ , \new_Sorter100|5660_ ,
    \new_Sorter100|5661_ , \new_Sorter100|5662_ , \new_Sorter100|5663_ ,
    \new_Sorter100|5664_ , \new_Sorter100|5665_ , \new_Sorter100|5666_ ,
    \new_Sorter100|5667_ , \new_Sorter100|5668_ , \new_Sorter100|5669_ ,
    \new_Sorter100|5670_ , \new_Sorter100|5671_ , \new_Sorter100|5672_ ,
    \new_Sorter100|5673_ , \new_Sorter100|5674_ , \new_Sorter100|5675_ ,
    \new_Sorter100|5676_ , \new_Sorter100|5677_ , \new_Sorter100|5678_ ,
    \new_Sorter100|5679_ , \new_Sorter100|5680_ , \new_Sorter100|5681_ ,
    \new_Sorter100|5682_ , \new_Sorter100|5683_ , \new_Sorter100|5684_ ,
    \new_Sorter100|5685_ , \new_Sorter100|5686_ , \new_Sorter100|5687_ ,
    \new_Sorter100|5688_ , \new_Sorter100|5689_ , \new_Sorter100|5690_ ,
    \new_Sorter100|5691_ , \new_Sorter100|5692_ , \new_Sorter100|5693_ ,
    \new_Sorter100|5694_ , \new_Sorter100|5695_ , \new_Sorter100|5696_ ,
    \new_Sorter100|5697_ , \new_Sorter100|5698_ , \new_Sorter100|5699_ ,
    \new_Sorter100|5700_ , \new_Sorter100|5799_ , \new_Sorter100|5701_ ,
    \new_Sorter100|5702_ , \new_Sorter100|5703_ , \new_Sorter100|5704_ ,
    \new_Sorter100|5705_ , \new_Sorter100|5706_ , \new_Sorter100|5707_ ,
    \new_Sorter100|5708_ , \new_Sorter100|5709_ , \new_Sorter100|5710_ ,
    \new_Sorter100|5711_ , \new_Sorter100|5712_ , \new_Sorter100|5713_ ,
    \new_Sorter100|5714_ , \new_Sorter100|5715_ , \new_Sorter100|5716_ ,
    \new_Sorter100|5717_ , \new_Sorter100|5718_ , \new_Sorter100|5719_ ,
    \new_Sorter100|5720_ , \new_Sorter100|5721_ , \new_Sorter100|5722_ ,
    \new_Sorter100|5723_ , \new_Sorter100|5724_ , \new_Sorter100|5725_ ,
    \new_Sorter100|5726_ , \new_Sorter100|5727_ , \new_Sorter100|5728_ ,
    \new_Sorter100|5729_ , \new_Sorter100|5730_ , \new_Sorter100|5731_ ,
    \new_Sorter100|5732_ , \new_Sorter100|5733_ , \new_Sorter100|5734_ ,
    \new_Sorter100|5735_ , \new_Sorter100|5736_ , \new_Sorter100|5737_ ,
    \new_Sorter100|5738_ , \new_Sorter100|5739_ , \new_Sorter100|5740_ ,
    \new_Sorter100|5741_ , \new_Sorter100|5742_ , \new_Sorter100|5743_ ,
    \new_Sorter100|5744_ , \new_Sorter100|5745_ , \new_Sorter100|5746_ ,
    \new_Sorter100|5747_ , \new_Sorter100|5748_ , \new_Sorter100|5749_ ,
    \new_Sorter100|5750_ , \new_Sorter100|5751_ , \new_Sorter100|5752_ ,
    \new_Sorter100|5753_ , \new_Sorter100|5754_ , \new_Sorter100|5755_ ,
    \new_Sorter100|5756_ , \new_Sorter100|5757_ , \new_Sorter100|5758_ ,
    \new_Sorter100|5759_ , \new_Sorter100|5760_ , \new_Sorter100|5761_ ,
    \new_Sorter100|5762_ , \new_Sorter100|5763_ , \new_Sorter100|5764_ ,
    \new_Sorter100|5765_ , \new_Sorter100|5766_ , \new_Sorter100|5767_ ,
    \new_Sorter100|5768_ , \new_Sorter100|5769_ , \new_Sorter100|5770_ ,
    \new_Sorter100|5771_ , \new_Sorter100|5772_ , \new_Sorter100|5773_ ,
    \new_Sorter100|5774_ , \new_Sorter100|5775_ , \new_Sorter100|5776_ ,
    \new_Sorter100|5777_ , \new_Sorter100|5778_ , \new_Sorter100|5779_ ,
    \new_Sorter100|5780_ , \new_Sorter100|5781_ , \new_Sorter100|5782_ ,
    \new_Sorter100|5783_ , \new_Sorter100|5784_ , \new_Sorter100|5785_ ,
    \new_Sorter100|5786_ , \new_Sorter100|5787_ , \new_Sorter100|5788_ ,
    \new_Sorter100|5789_ , \new_Sorter100|5790_ , \new_Sorter100|5791_ ,
    \new_Sorter100|5792_ , \new_Sorter100|5793_ , \new_Sorter100|5794_ ,
    \new_Sorter100|5795_ , \new_Sorter100|5796_ , \new_Sorter100|5797_ ,
    \new_Sorter100|5798_ , \new_Sorter100|5800_ , \new_Sorter100|5801_ ,
    \new_Sorter100|5802_ , \new_Sorter100|5803_ , \new_Sorter100|5804_ ,
    \new_Sorter100|5805_ , \new_Sorter100|5806_ , \new_Sorter100|5807_ ,
    \new_Sorter100|5808_ , \new_Sorter100|5809_ , \new_Sorter100|5810_ ,
    \new_Sorter100|5811_ , \new_Sorter100|5812_ , \new_Sorter100|5813_ ,
    \new_Sorter100|5814_ , \new_Sorter100|5815_ , \new_Sorter100|5816_ ,
    \new_Sorter100|5817_ , \new_Sorter100|5818_ , \new_Sorter100|5819_ ,
    \new_Sorter100|5820_ , \new_Sorter100|5821_ , \new_Sorter100|5822_ ,
    \new_Sorter100|5823_ , \new_Sorter100|5824_ , \new_Sorter100|5825_ ,
    \new_Sorter100|5826_ , \new_Sorter100|5827_ , \new_Sorter100|5828_ ,
    \new_Sorter100|5829_ , \new_Sorter100|5830_ , \new_Sorter100|5831_ ,
    \new_Sorter100|5832_ , \new_Sorter100|5833_ , \new_Sorter100|5834_ ,
    \new_Sorter100|5835_ , \new_Sorter100|5836_ , \new_Sorter100|5837_ ,
    \new_Sorter100|5838_ , \new_Sorter100|5839_ , \new_Sorter100|5840_ ,
    \new_Sorter100|5841_ , \new_Sorter100|5842_ , \new_Sorter100|5843_ ,
    \new_Sorter100|5844_ , \new_Sorter100|5845_ , \new_Sorter100|5846_ ,
    \new_Sorter100|5847_ , \new_Sorter100|5848_ , \new_Sorter100|5849_ ,
    \new_Sorter100|5850_ , \new_Sorter100|5851_ , \new_Sorter100|5852_ ,
    \new_Sorter100|5853_ , \new_Sorter100|5854_ , \new_Sorter100|5855_ ,
    \new_Sorter100|5856_ , \new_Sorter100|5857_ , \new_Sorter100|5858_ ,
    \new_Sorter100|5859_ , \new_Sorter100|5860_ , \new_Sorter100|5861_ ,
    \new_Sorter100|5862_ , \new_Sorter100|5863_ , \new_Sorter100|5864_ ,
    \new_Sorter100|5865_ , \new_Sorter100|5866_ , \new_Sorter100|5867_ ,
    \new_Sorter100|5868_ , \new_Sorter100|5869_ , \new_Sorter100|5870_ ,
    \new_Sorter100|5871_ , \new_Sorter100|5872_ , \new_Sorter100|5873_ ,
    \new_Sorter100|5874_ , \new_Sorter100|5875_ , \new_Sorter100|5876_ ,
    \new_Sorter100|5877_ , \new_Sorter100|5878_ , \new_Sorter100|5879_ ,
    \new_Sorter100|5880_ , \new_Sorter100|5881_ , \new_Sorter100|5882_ ,
    \new_Sorter100|5883_ , \new_Sorter100|5884_ , \new_Sorter100|5885_ ,
    \new_Sorter100|5886_ , \new_Sorter100|5887_ , \new_Sorter100|5888_ ,
    \new_Sorter100|5889_ , \new_Sorter100|5890_ , \new_Sorter100|5891_ ,
    \new_Sorter100|5892_ , \new_Sorter100|5893_ , \new_Sorter100|5894_ ,
    \new_Sorter100|5895_ , \new_Sorter100|5896_ , \new_Sorter100|5897_ ,
    \new_Sorter100|5898_ , \new_Sorter100|5899_ , \new_Sorter100|5900_ ,
    \new_Sorter100|5999_ , \new_Sorter100|5901_ , \new_Sorter100|5902_ ,
    \new_Sorter100|5903_ , \new_Sorter100|5904_ , \new_Sorter100|5905_ ,
    \new_Sorter100|5906_ , \new_Sorter100|5907_ , \new_Sorter100|5908_ ,
    \new_Sorter100|5909_ , \new_Sorter100|5910_ , \new_Sorter100|5911_ ,
    \new_Sorter100|5912_ , \new_Sorter100|5913_ , \new_Sorter100|5914_ ,
    \new_Sorter100|5915_ , \new_Sorter100|5916_ , \new_Sorter100|5917_ ,
    \new_Sorter100|5918_ , \new_Sorter100|5919_ , \new_Sorter100|5920_ ,
    \new_Sorter100|5921_ , \new_Sorter100|5922_ , \new_Sorter100|5923_ ,
    \new_Sorter100|5924_ , \new_Sorter100|5925_ , \new_Sorter100|5926_ ,
    \new_Sorter100|5927_ , \new_Sorter100|5928_ , \new_Sorter100|5929_ ,
    \new_Sorter100|5930_ , \new_Sorter100|5931_ , \new_Sorter100|5932_ ,
    \new_Sorter100|5933_ , \new_Sorter100|5934_ , \new_Sorter100|5935_ ,
    \new_Sorter100|5936_ , \new_Sorter100|5937_ , \new_Sorter100|5938_ ,
    \new_Sorter100|5939_ , \new_Sorter100|5940_ , \new_Sorter100|5941_ ,
    \new_Sorter100|5942_ , \new_Sorter100|5943_ , \new_Sorter100|5944_ ,
    \new_Sorter100|5945_ , \new_Sorter100|5946_ , \new_Sorter100|5947_ ,
    \new_Sorter100|5948_ , \new_Sorter100|5949_ , \new_Sorter100|5950_ ,
    \new_Sorter100|5951_ , \new_Sorter100|5952_ , \new_Sorter100|5953_ ,
    \new_Sorter100|5954_ , \new_Sorter100|5955_ , \new_Sorter100|5956_ ,
    \new_Sorter100|5957_ , \new_Sorter100|5958_ , \new_Sorter100|5959_ ,
    \new_Sorter100|5960_ , \new_Sorter100|5961_ , \new_Sorter100|5962_ ,
    \new_Sorter100|5963_ , \new_Sorter100|5964_ , \new_Sorter100|5965_ ,
    \new_Sorter100|5966_ , \new_Sorter100|5967_ , \new_Sorter100|5968_ ,
    \new_Sorter100|5969_ , \new_Sorter100|5970_ , \new_Sorter100|5971_ ,
    \new_Sorter100|5972_ , \new_Sorter100|5973_ , \new_Sorter100|5974_ ,
    \new_Sorter100|5975_ , \new_Sorter100|5976_ , \new_Sorter100|5977_ ,
    \new_Sorter100|5978_ , \new_Sorter100|5979_ , \new_Sorter100|5980_ ,
    \new_Sorter100|5981_ , \new_Sorter100|5982_ , \new_Sorter100|5983_ ,
    \new_Sorter100|5984_ , \new_Sorter100|5985_ , \new_Sorter100|5986_ ,
    \new_Sorter100|5987_ , \new_Sorter100|5988_ , \new_Sorter100|5989_ ,
    \new_Sorter100|5990_ , \new_Sorter100|5991_ , \new_Sorter100|5992_ ,
    \new_Sorter100|5993_ , \new_Sorter100|5994_ , \new_Sorter100|5995_ ,
    \new_Sorter100|5996_ , \new_Sorter100|5997_ , \new_Sorter100|5998_ ,
    \new_Sorter100|6000_ , \new_Sorter100|6001_ , \new_Sorter100|6002_ ,
    \new_Sorter100|6003_ , \new_Sorter100|6004_ , \new_Sorter100|6005_ ,
    \new_Sorter100|6006_ , \new_Sorter100|6007_ , \new_Sorter100|6008_ ,
    \new_Sorter100|6009_ , \new_Sorter100|6010_ , \new_Sorter100|6011_ ,
    \new_Sorter100|6012_ , \new_Sorter100|6013_ , \new_Sorter100|6014_ ,
    \new_Sorter100|6015_ , \new_Sorter100|6016_ , \new_Sorter100|6017_ ,
    \new_Sorter100|6018_ , \new_Sorter100|6019_ , \new_Sorter100|6020_ ,
    \new_Sorter100|6021_ , \new_Sorter100|6022_ , \new_Sorter100|6023_ ,
    \new_Sorter100|6024_ , \new_Sorter100|6025_ , \new_Sorter100|6026_ ,
    \new_Sorter100|6027_ , \new_Sorter100|6028_ , \new_Sorter100|6029_ ,
    \new_Sorter100|6030_ , \new_Sorter100|6031_ , \new_Sorter100|6032_ ,
    \new_Sorter100|6033_ , \new_Sorter100|6034_ , \new_Sorter100|6035_ ,
    \new_Sorter100|6036_ , \new_Sorter100|6037_ , \new_Sorter100|6038_ ,
    \new_Sorter100|6039_ , \new_Sorter100|6040_ , \new_Sorter100|6041_ ,
    \new_Sorter100|6042_ , \new_Sorter100|6043_ , \new_Sorter100|6044_ ,
    \new_Sorter100|6045_ , \new_Sorter100|6046_ , \new_Sorter100|6047_ ,
    \new_Sorter100|6048_ , \new_Sorter100|6049_ , \new_Sorter100|6050_ ,
    \new_Sorter100|6051_ , \new_Sorter100|6052_ , \new_Sorter100|6053_ ,
    \new_Sorter100|6054_ , \new_Sorter100|6055_ , \new_Sorter100|6056_ ,
    \new_Sorter100|6057_ , \new_Sorter100|6058_ , \new_Sorter100|6059_ ,
    \new_Sorter100|6060_ , \new_Sorter100|6061_ , \new_Sorter100|6062_ ,
    \new_Sorter100|6063_ , \new_Sorter100|6064_ , \new_Sorter100|6065_ ,
    \new_Sorter100|6066_ , \new_Sorter100|6067_ , \new_Sorter100|6068_ ,
    \new_Sorter100|6069_ , \new_Sorter100|6070_ , \new_Sorter100|6071_ ,
    \new_Sorter100|6072_ , \new_Sorter100|6073_ , \new_Sorter100|6074_ ,
    \new_Sorter100|6075_ , \new_Sorter100|6076_ , \new_Sorter100|6077_ ,
    \new_Sorter100|6078_ , \new_Sorter100|6079_ , \new_Sorter100|6080_ ,
    \new_Sorter100|6081_ , \new_Sorter100|6082_ , \new_Sorter100|6083_ ,
    \new_Sorter100|6084_ , \new_Sorter100|6085_ , \new_Sorter100|6086_ ,
    \new_Sorter100|6087_ , \new_Sorter100|6088_ , \new_Sorter100|6089_ ,
    \new_Sorter100|6090_ , \new_Sorter100|6091_ , \new_Sorter100|6092_ ,
    \new_Sorter100|6093_ , \new_Sorter100|6094_ , \new_Sorter100|6095_ ,
    \new_Sorter100|6096_ , \new_Sorter100|6097_ , \new_Sorter100|6098_ ,
    \new_Sorter100|6099_ , \new_Sorter100|6100_ , \new_Sorter100|6199_ ,
    \new_Sorter100|6101_ , \new_Sorter100|6102_ , \new_Sorter100|6103_ ,
    \new_Sorter100|6104_ , \new_Sorter100|6105_ , \new_Sorter100|6106_ ,
    \new_Sorter100|6107_ , \new_Sorter100|6108_ , \new_Sorter100|6109_ ,
    \new_Sorter100|6110_ , \new_Sorter100|6111_ , \new_Sorter100|6112_ ,
    \new_Sorter100|6113_ , \new_Sorter100|6114_ , \new_Sorter100|6115_ ,
    \new_Sorter100|6116_ , \new_Sorter100|6117_ , \new_Sorter100|6118_ ,
    \new_Sorter100|6119_ , \new_Sorter100|6120_ , \new_Sorter100|6121_ ,
    \new_Sorter100|6122_ , \new_Sorter100|6123_ , \new_Sorter100|6124_ ,
    \new_Sorter100|6125_ , \new_Sorter100|6126_ , \new_Sorter100|6127_ ,
    \new_Sorter100|6128_ , \new_Sorter100|6129_ , \new_Sorter100|6130_ ,
    \new_Sorter100|6131_ , \new_Sorter100|6132_ , \new_Sorter100|6133_ ,
    \new_Sorter100|6134_ , \new_Sorter100|6135_ , \new_Sorter100|6136_ ,
    \new_Sorter100|6137_ , \new_Sorter100|6138_ , \new_Sorter100|6139_ ,
    \new_Sorter100|6140_ , \new_Sorter100|6141_ , \new_Sorter100|6142_ ,
    \new_Sorter100|6143_ , \new_Sorter100|6144_ , \new_Sorter100|6145_ ,
    \new_Sorter100|6146_ , \new_Sorter100|6147_ , \new_Sorter100|6148_ ,
    \new_Sorter100|6149_ , \new_Sorter100|6150_ , \new_Sorter100|6151_ ,
    \new_Sorter100|6152_ , \new_Sorter100|6153_ , \new_Sorter100|6154_ ,
    \new_Sorter100|6155_ , \new_Sorter100|6156_ , \new_Sorter100|6157_ ,
    \new_Sorter100|6158_ , \new_Sorter100|6159_ , \new_Sorter100|6160_ ,
    \new_Sorter100|6161_ , \new_Sorter100|6162_ , \new_Sorter100|6163_ ,
    \new_Sorter100|6164_ , \new_Sorter100|6165_ , \new_Sorter100|6166_ ,
    \new_Sorter100|6167_ , \new_Sorter100|6168_ , \new_Sorter100|6169_ ,
    \new_Sorter100|6170_ , \new_Sorter100|6171_ , \new_Sorter100|6172_ ,
    \new_Sorter100|6173_ , \new_Sorter100|6174_ , \new_Sorter100|6175_ ,
    \new_Sorter100|6176_ , \new_Sorter100|6177_ , \new_Sorter100|6178_ ,
    \new_Sorter100|6179_ , \new_Sorter100|6180_ , \new_Sorter100|6181_ ,
    \new_Sorter100|6182_ , \new_Sorter100|6183_ , \new_Sorter100|6184_ ,
    \new_Sorter100|6185_ , \new_Sorter100|6186_ , \new_Sorter100|6187_ ,
    \new_Sorter100|6188_ , \new_Sorter100|6189_ , \new_Sorter100|6190_ ,
    \new_Sorter100|6191_ , \new_Sorter100|6192_ , \new_Sorter100|6193_ ,
    \new_Sorter100|6194_ , \new_Sorter100|6195_ , \new_Sorter100|6196_ ,
    \new_Sorter100|6197_ , \new_Sorter100|6198_ , \new_Sorter100|6200_ ,
    \new_Sorter100|6201_ , \new_Sorter100|6202_ , \new_Sorter100|6203_ ,
    \new_Sorter100|6204_ , \new_Sorter100|6205_ , \new_Sorter100|6206_ ,
    \new_Sorter100|6207_ , \new_Sorter100|6208_ , \new_Sorter100|6209_ ,
    \new_Sorter100|6210_ , \new_Sorter100|6211_ , \new_Sorter100|6212_ ,
    \new_Sorter100|6213_ , \new_Sorter100|6214_ , \new_Sorter100|6215_ ,
    \new_Sorter100|6216_ , \new_Sorter100|6217_ , \new_Sorter100|6218_ ,
    \new_Sorter100|6219_ , \new_Sorter100|6220_ , \new_Sorter100|6221_ ,
    \new_Sorter100|6222_ , \new_Sorter100|6223_ , \new_Sorter100|6224_ ,
    \new_Sorter100|6225_ , \new_Sorter100|6226_ , \new_Sorter100|6227_ ,
    \new_Sorter100|6228_ , \new_Sorter100|6229_ , \new_Sorter100|6230_ ,
    \new_Sorter100|6231_ , \new_Sorter100|6232_ , \new_Sorter100|6233_ ,
    \new_Sorter100|6234_ , \new_Sorter100|6235_ , \new_Sorter100|6236_ ,
    \new_Sorter100|6237_ , \new_Sorter100|6238_ , \new_Sorter100|6239_ ,
    \new_Sorter100|6240_ , \new_Sorter100|6241_ , \new_Sorter100|6242_ ,
    \new_Sorter100|6243_ , \new_Sorter100|6244_ , \new_Sorter100|6245_ ,
    \new_Sorter100|6246_ , \new_Sorter100|6247_ , \new_Sorter100|6248_ ,
    \new_Sorter100|6249_ , \new_Sorter100|6250_ , \new_Sorter100|6251_ ,
    \new_Sorter100|6252_ , \new_Sorter100|6253_ , \new_Sorter100|6254_ ,
    \new_Sorter100|6255_ , \new_Sorter100|6256_ , \new_Sorter100|6257_ ,
    \new_Sorter100|6258_ , \new_Sorter100|6259_ , \new_Sorter100|6260_ ,
    \new_Sorter100|6261_ , \new_Sorter100|6262_ , \new_Sorter100|6263_ ,
    \new_Sorter100|6264_ , \new_Sorter100|6265_ , \new_Sorter100|6266_ ,
    \new_Sorter100|6267_ , \new_Sorter100|6268_ , \new_Sorter100|6269_ ,
    \new_Sorter100|6270_ , \new_Sorter100|6271_ , \new_Sorter100|6272_ ,
    \new_Sorter100|6273_ , \new_Sorter100|6274_ , \new_Sorter100|6275_ ,
    \new_Sorter100|6276_ , \new_Sorter100|6277_ , \new_Sorter100|6278_ ,
    \new_Sorter100|6279_ , \new_Sorter100|6280_ , \new_Sorter100|6281_ ,
    \new_Sorter100|6282_ , \new_Sorter100|6283_ , \new_Sorter100|6284_ ,
    \new_Sorter100|6285_ , \new_Sorter100|6286_ , \new_Sorter100|6287_ ,
    \new_Sorter100|6288_ , \new_Sorter100|6289_ , \new_Sorter100|6290_ ,
    \new_Sorter100|6291_ , \new_Sorter100|6292_ , \new_Sorter100|6293_ ,
    \new_Sorter100|6294_ , \new_Sorter100|6295_ , \new_Sorter100|6296_ ,
    \new_Sorter100|6297_ , \new_Sorter100|6298_ , \new_Sorter100|6299_ ,
    \new_Sorter100|6300_ , \new_Sorter100|6399_ , \new_Sorter100|6301_ ,
    \new_Sorter100|6302_ , \new_Sorter100|6303_ , \new_Sorter100|6304_ ,
    \new_Sorter100|6305_ , \new_Sorter100|6306_ , \new_Sorter100|6307_ ,
    \new_Sorter100|6308_ , \new_Sorter100|6309_ , \new_Sorter100|6310_ ,
    \new_Sorter100|6311_ , \new_Sorter100|6312_ , \new_Sorter100|6313_ ,
    \new_Sorter100|6314_ , \new_Sorter100|6315_ , \new_Sorter100|6316_ ,
    \new_Sorter100|6317_ , \new_Sorter100|6318_ , \new_Sorter100|6319_ ,
    \new_Sorter100|6320_ , \new_Sorter100|6321_ , \new_Sorter100|6322_ ,
    \new_Sorter100|6323_ , \new_Sorter100|6324_ , \new_Sorter100|6325_ ,
    \new_Sorter100|6326_ , \new_Sorter100|6327_ , \new_Sorter100|6328_ ,
    \new_Sorter100|6329_ , \new_Sorter100|6330_ , \new_Sorter100|6331_ ,
    \new_Sorter100|6332_ , \new_Sorter100|6333_ , \new_Sorter100|6334_ ,
    \new_Sorter100|6335_ , \new_Sorter100|6336_ , \new_Sorter100|6337_ ,
    \new_Sorter100|6338_ , \new_Sorter100|6339_ , \new_Sorter100|6340_ ,
    \new_Sorter100|6341_ , \new_Sorter100|6342_ , \new_Sorter100|6343_ ,
    \new_Sorter100|6344_ , \new_Sorter100|6345_ , \new_Sorter100|6346_ ,
    \new_Sorter100|6347_ , \new_Sorter100|6348_ , \new_Sorter100|6349_ ,
    \new_Sorter100|6350_ , \new_Sorter100|6351_ , \new_Sorter100|6352_ ,
    \new_Sorter100|6353_ , \new_Sorter100|6354_ , \new_Sorter100|6355_ ,
    \new_Sorter100|6356_ , \new_Sorter100|6357_ , \new_Sorter100|6358_ ,
    \new_Sorter100|6359_ , \new_Sorter100|6360_ , \new_Sorter100|6361_ ,
    \new_Sorter100|6362_ , \new_Sorter100|6363_ , \new_Sorter100|6364_ ,
    \new_Sorter100|6365_ , \new_Sorter100|6366_ , \new_Sorter100|6367_ ,
    \new_Sorter100|6368_ , \new_Sorter100|6369_ , \new_Sorter100|6370_ ,
    \new_Sorter100|6371_ , \new_Sorter100|6372_ , \new_Sorter100|6373_ ,
    \new_Sorter100|6374_ , \new_Sorter100|6375_ , \new_Sorter100|6376_ ,
    \new_Sorter100|6377_ , \new_Sorter100|6378_ , \new_Sorter100|6379_ ,
    \new_Sorter100|6380_ , \new_Sorter100|6381_ , \new_Sorter100|6382_ ,
    \new_Sorter100|6383_ , \new_Sorter100|6384_ , \new_Sorter100|6385_ ,
    \new_Sorter100|6386_ , \new_Sorter100|6387_ , \new_Sorter100|6388_ ,
    \new_Sorter100|6389_ , \new_Sorter100|6390_ , \new_Sorter100|6391_ ,
    \new_Sorter100|6392_ , \new_Sorter100|6393_ , \new_Sorter100|6394_ ,
    \new_Sorter100|6395_ , \new_Sorter100|6396_ , \new_Sorter100|6397_ ,
    \new_Sorter100|6398_ , \new_Sorter100|6400_ , \new_Sorter100|6401_ ,
    \new_Sorter100|6402_ , \new_Sorter100|6403_ , \new_Sorter100|6404_ ,
    \new_Sorter100|6405_ , \new_Sorter100|6406_ , \new_Sorter100|6407_ ,
    \new_Sorter100|6408_ , \new_Sorter100|6409_ , \new_Sorter100|6410_ ,
    \new_Sorter100|6411_ , \new_Sorter100|6412_ , \new_Sorter100|6413_ ,
    \new_Sorter100|6414_ , \new_Sorter100|6415_ , \new_Sorter100|6416_ ,
    \new_Sorter100|6417_ , \new_Sorter100|6418_ , \new_Sorter100|6419_ ,
    \new_Sorter100|6420_ , \new_Sorter100|6421_ , \new_Sorter100|6422_ ,
    \new_Sorter100|6423_ , \new_Sorter100|6424_ , \new_Sorter100|6425_ ,
    \new_Sorter100|6426_ , \new_Sorter100|6427_ , \new_Sorter100|6428_ ,
    \new_Sorter100|6429_ , \new_Sorter100|6430_ , \new_Sorter100|6431_ ,
    \new_Sorter100|6432_ , \new_Sorter100|6433_ , \new_Sorter100|6434_ ,
    \new_Sorter100|6435_ , \new_Sorter100|6436_ , \new_Sorter100|6437_ ,
    \new_Sorter100|6438_ , \new_Sorter100|6439_ , \new_Sorter100|6440_ ,
    \new_Sorter100|6441_ , \new_Sorter100|6442_ , \new_Sorter100|6443_ ,
    \new_Sorter100|6444_ , \new_Sorter100|6445_ , \new_Sorter100|6446_ ,
    \new_Sorter100|6447_ , \new_Sorter100|6448_ , \new_Sorter100|6449_ ,
    \new_Sorter100|6450_ , \new_Sorter100|6451_ , \new_Sorter100|6452_ ,
    \new_Sorter100|6453_ , \new_Sorter100|6454_ , \new_Sorter100|6455_ ,
    \new_Sorter100|6456_ , \new_Sorter100|6457_ , \new_Sorter100|6458_ ,
    \new_Sorter100|6459_ , \new_Sorter100|6460_ , \new_Sorter100|6461_ ,
    \new_Sorter100|6462_ , \new_Sorter100|6463_ , \new_Sorter100|6464_ ,
    \new_Sorter100|6465_ , \new_Sorter100|6466_ , \new_Sorter100|6467_ ,
    \new_Sorter100|6468_ , \new_Sorter100|6469_ , \new_Sorter100|6470_ ,
    \new_Sorter100|6471_ , \new_Sorter100|6472_ , \new_Sorter100|6473_ ,
    \new_Sorter100|6474_ , \new_Sorter100|6475_ , \new_Sorter100|6476_ ,
    \new_Sorter100|6477_ , \new_Sorter100|6478_ , \new_Sorter100|6479_ ,
    \new_Sorter100|6480_ , \new_Sorter100|6481_ , \new_Sorter100|6482_ ,
    \new_Sorter100|6483_ , \new_Sorter100|6484_ , \new_Sorter100|6485_ ,
    \new_Sorter100|6486_ , \new_Sorter100|6487_ , \new_Sorter100|6488_ ,
    \new_Sorter100|6489_ , \new_Sorter100|6490_ , \new_Sorter100|6491_ ,
    \new_Sorter100|6492_ , \new_Sorter100|6493_ , \new_Sorter100|6494_ ,
    \new_Sorter100|6495_ , \new_Sorter100|6496_ , \new_Sorter100|6497_ ,
    \new_Sorter100|6498_ , \new_Sorter100|6499_ , \new_Sorter100|6500_ ,
    \new_Sorter100|6599_ , \new_Sorter100|6501_ , \new_Sorter100|6502_ ,
    \new_Sorter100|6503_ , \new_Sorter100|6504_ , \new_Sorter100|6505_ ,
    \new_Sorter100|6506_ , \new_Sorter100|6507_ , \new_Sorter100|6508_ ,
    \new_Sorter100|6509_ , \new_Sorter100|6510_ , \new_Sorter100|6511_ ,
    \new_Sorter100|6512_ , \new_Sorter100|6513_ , \new_Sorter100|6514_ ,
    \new_Sorter100|6515_ , \new_Sorter100|6516_ , \new_Sorter100|6517_ ,
    \new_Sorter100|6518_ , \new_Sorter100|6519_ , \new_Sorter100|6520_ ,
    \new_Sorter100|6521_ , \new_Sorter100|6522_ , \new_Sorter100|6523_ ,
    \new_Sorter100|6524_ , \new_Sorter100|6525_ , \new_Sorter100|6526_ ,
    \new_Sorter100|6527_ , \new_Sorter100|6528_ , \new_Sorter100|6529_ ,
    \new_Sorter100|6530_ , \new_Sorter100|6531_ , \new_Sorter100|6532_ ,
    \new_Sorter100|6533_ , \new_Sorter100|6534_ , \new_Sorter100|6535_ ,
    \new_Sorter100|6536_ , \new_Sorter100|6537_ , \new_Sorter100|6538_ ,
    \new_Sorter100|6539_ , \new_Sorter100|6540_ , \new_Sorter100|6541_ ,
    \new_Sorter100|6542_ , \new_Sorter100|6543_ , \new_Sorter100|6544_ ,
    \new_Sorter100|6545_ , \new_Sorter100|6546_ , \new_Sorter100|6547_ ,
    \new_Sorter100|6548_ , \new_Sorter100|6549_ , \new_Sorter100|6550_ ,
    \new_Sorter100|6551_ , \new_Sorter100|6552_ , \new_Sorter100|6553_ ,
    \new_Sorter100|6554_ , \new_Sorter100|6555_ , \new_Sorter100|6556_ ,
    \new_Sorter100|6557_ , \new_Sorter100|6558_ , \new_Sorter100|6559_ ,
    \new_Sorter100|6560_ , \new_Sorter100|6561_ , \new_Sorter100|6562_ ,
    \new_Sorter100|6563_ , \new_Sorter100|6564_ , \new_Sorter100|6565_ ,
    \new_Sorter100|6566_ , \new_Sorter100|6567_ , \new_Sorter100|6568_ ,
    \new_Sorter100|6569_ , \new_Sorter100|6570_ , \new_Sorter100|6571_ ,
    \new_Sorter100|6572_ , \new_Sorter100|6573_ , \new_Sorter100|6574_ ,
    \new_Sorter100|6575_ , \new_Sorter100|6576_ , \new_Sorter100|6577_ ,
    \new_Sorter100|6578_ , \new_Sorter100|6579_ , \new_Sorter100|6580_ ,
    \new_Sorter100|6581_ , \new_Sorter100|6582_ , \new_Sorter100|6583_ ,
    \new_Sorter100|6584_ , \new_Sorter100|6585_ , \new_Sorter100|6586_ ,
    \new_Sorter100|6587_ , \new_Sorter100|6588_ , \new_Sorter100|6589_ ,
    \new_Sorter100|6590_ , \new_Sorter100|6591_ , \new_Sorter100|6592_ ,
    \new_Sorter100|6593_ , \new_Sorter100|6594_ , \new_Sorter100|6595_ ,
    \new_Sorter100|6596_ , \new_Sorter100|6597_ , \new_Sorter100|6598_ ,
    \new_Sorter100|6600_ , \new_Sorter100|6601_ , \new_Sorter100|6602_ ,
    \new_Sorter100|6603_ , \new_Sorter100|6604_ , \new_Sorter100|6605_ ,
    \new_Sorter100|6606_ , \new_Sorter100|6607_ , \new_Sorter100|6608_ ,
    \new_Sorter100|6609_ , \new_Sorter100|6610_ , \new_Sorter100|6611_ ,
    \new_Sorter100|6612_ , \new_Sorter100|6613_ , \new_Sorter100|6614_ ,
    \new_Sorter100|6615_ , \new_Sorter100|6616_ , \new_Sorter100|6617_ ,
    \new_Sorter100|6618_ , \new_Sorter100|6619_ , \new_Sorter100|6620_ ,
    \new_Sorter100|6621_ , \new_Sorter100|6622_ , \new_Sorter100|6623_ ,
    \new_Sorter100|6624_ , \new_Sorter100|6625_ , \new_Sorter100|6626_ ,
    \new_Sorter100|6627_ , \new_Sorter100|6628_ , \new_Sorter100|6629_ ,
    \new_Sorter100|6630_ , \new_Sorter100|6631_ , \new_Sorter100|6632_ ,
    \new_Sorter100|6633_ , \new_Sorter100|6634_ , \new_Sorter100|6635_ ,
    \new_Sorter100|6636_ , \new_Sorter100|6637_ , \new_Sorter100|6638_ ,
    \new_Sorter100|6639_ , \new_Sorter100|6640_ , \new_Sorter100|6641_ ,
    \new_Sorter100|6642_ , \new_Sorter100|6643_ , \new_Sorter100|6644_ ,
    \new_Sorter100|6645_ , \new_Sorter100|6646_ , \new_Sorter100|6647_ ,
    \new_Sorter100|6648_ , \new_Sorter100|6649_ , \new_Sorter100|6650_ ,
    \new_Sorter100|6651_ , \new_Sorter100|6652_ , \new_Sorter100|6653_ ,
    \new_Sorter100|6654_ , \new_Sorter100|6655_ , \new_Sorter100|6656_ ,
    \new_Sorter100|6657_ , \new_Sorter100|6658_ , \new_Sorter100|6659_ ,
    \new_Sorter100|6660_ , \new_Sorter100|6661_ , \new_Sorter100|6662_ ,
    \new_Sorter100|6663_ , \new_Sorter100|6664_ , \new_Sorter100|6665_ ,
    \new_Sorter100|6666_ , \new_Sorter100|6667_ , \new_Sorter100|6668_ ,
    \new_Sorter100|6669_ , \new_Sorter100|6670_ , \new_Sorter100|6671_ ,
    \new_Sorter100|6672_ , \new_Sorter100|6673_ , \new_Sorter100|6674_ ,
    \new_Sorter100|6675_ , \new_Sorter100|6676_ , \new_Sorter100|6677_ ,
    \new_Sorter100|6678_ , \new_Sorter100|6679_ , \new_Sorter100|6680_ ,
    \new_Sorter100|6681_ , \new_Sorter100|6682_ , \new_Sorter100|6683_ ,
    \new_Sorter100|6684_ , \new_Sorter100|6685_ , \new_Sorter100|6686_ ,
    \new_Sorter100|6687_ , \new_Sorter100|6688_ , \new_Sorter100|6689_ ,
    \new_Sorter100|6690_ , \new_Sorter100|6691_ , \new_Sorter100|6692_ ,
    \new_Sorter100|6693_ , \new_Sorter100|6694_ , \new_Sorter100|6695_ ,
    \new_Sorter100|6696_ , \new_Sorter100|6697_ , \new_Sorter100|6698_ ,
    \new_Sorter100|6699_ , \new_Sorter100|6700_ , \new_Sorter100|6799_ ,
    \new_Sorter100|6701_ , \new_Sorter100|6702_ , \new_Sorter100|6703_ ,
    \new_Sorter100|6704_ , \new_Sorter100|6705_ , \new_Sorter100|6706_ ,
    \new_Sorter100|6707_ , \new_Sorter100|6708_ , \new_Sorter100|6709_ ,
    \new_Sorter100|6710_ , \new_Sorter100|6711_ , \new_Sorter100|6712_ ,
    \new_Sorter100|6713_ , \new_Sorter100|6714_ , \new_Sorter100|6715_ ,
    \new_Sorter100|6716_ , \new_Sorter100|6717_ , \new_Sorter100|6718_ ,
    \new_Sorter100|6719_ , \new_Sorter100|6720_ , \new_Sorter100|6721_ ,
    \new_Sorter100|6722_ , \new_Sorter100|6723_ , \new_Sorter100|6724_ ,
    \new_Sorter100|6725_ , \new_Sorter100|6726_ , \new_Sorter100|6727_ ,
    \new_Sorter100|6728_ , \new_Sorter100|6729_ , \new_Sorter100|6730_ ,
    \new_Sorter100|6731_ , \new_Sorter100|6732_ , \new_Sorter100|6733_ ,
    \new_Sorter100|6734_ , \new_Sorter100|6735_ , \new_Sorter100|6736_ ,
    \new_Sorter100|6737_ , \new_Sorter100|6738_ , \new_Sorter100|6739_ ,
    \new_Sorter100|6740_ , \new_Sorter100|6741_ , \new_Sorter100|6742_ ,
    \new_Sorter100|6743_ , \new_Sorter100|6744_ , \new_Sorter100|6745_ ,
    \new_Sorter100|6746_ , \new_Sorter100|6747_ , \new_Sorter100|6748_ ,
    \new_Sorter100|6749_ , \new_Sorter100|6750_ , \new_Sorter100|6751_ ,
    \new_Sorter100|6752_ , \new_Sorter100|6753_ , \new_Sorter100|6754_ ,
    \new_Sorter100|6755_ , \new_Sorter100|6756_ , \new_Sorter100|6757_ ,
    \new_Sorter100|6758_ , \new_Sorter100|6759_ , \new_Sorter100|6760_ ,
    \new_Sorter100|6761_ , \new_Sorter100|6762_ , \new_Sorter100|6763_ ,
    \new_Sorter100|6764_ , \new_Sorter100|6765_ , \new_Sorter100|6766_ ,
    \new_Sorter100|6767_ , \new_Sorter100|6768_ , \new_Sorter100|6769_ ,
    \new_Sorter100|6770_ , \new_Sorter100|6771_ , \new_Sorter100|6772_ ,
    \new_Sorter100|6773_ , \new_Sorter100|6774_ , \new_Sorter100|6775_ ,
    \new_Sorter100|6776_ , \new_Sorter100|6777_ , \new_Sorter100|6778_ ,
    \new_Sorter100|6779_ , \new_Sorter100|6780_ , \new_Sorter100|6781_ ,
    \new_Sorter100|6782_ , \new_Sorter100|6783_ , \new_Sorter100|6784_ ,
    \new_Sorter100|6785_ , \new_Sorter100|6786_ , \new_Sorter100|6787_ ,
    \new_Sorter100|6788_ , \new_Sorter100|6789_ , \new_Sorter100|6790_ ,
    \new_Sorter100|6791_ , \new_Sorter100|6792_ , \new_Sorter100|6793_ ,
    \new_Sorter100|6794_ , \new_Sorter100|6795_ , \new_Sorter100|6796_ ,
    \new_Sorter100|6797_ , \new_Sorter100|6798_ , \new_Sorter100|6800_ ,
    \new_Sorter100|6801_ , \new_Sorter100|6802_ , \new_Sorter100|6803_ ,
    \new_Sorter100|6804_ , \new_Sorter100|6805_ , \new_Sorter100|6806_ ,
    \new_Sorter100|6807_ , \new_Sorter100|6808_ , \new_Sorter100|6809_ ,
    \new_Sorter100|6810_ , \new_Sorter100|6811_ , \new_Sorter100|6812_ ,
    \new_Sorter100|6813_ , \new_Sorter100|6814_ , \new_Sorter100|6815_ ,
    \new_Sorter100|6816_ , \new_Sorter100|6817_ , \new_Sorter100|6818_ ,
    \new_Sorter100|6819_ , \new_Sorter100|6820_ , \new_Sorter100|6821_ ,
    \new_Sorter100|6822_ , \new_Sorter100|6823_ , \new_Sorter100|6824_ ,
    \new_Sorter100|6825_ , \new_Sorter100|6826_ , \new_Sorter100|6827_ ,
    \new_Sorter100|6828_ , \new_Sorter100|6829_ , \new_Sorter100|6830_ ,
    \new_Sorter100|6831_ , \new_Sorter100|6832_ , \new_Sorter100|6833_ ,
    \new_Sorter100|6834_ , \new_Sorter100|6835_ , \new_Sorter100|6836_ ,
    \new_Sorter100|6837_ , \new_Sorter100|6838_ , \new_Sorter100|6839_ ,
    \new_Sorter100|6840_ , \new_Sorter100|6841_ , \new_Sorter100|6842_ ,
    \new_Sorter100|6843_ , \new_Sorter100|6844_ , \new_Sorter100|6845_ ,
    \new_Sorter100|6846_ , \new_Sorter100|6847_ , \new_Sorter100|6848_ ,
    \new_Sorter100|6849_ , \new_Sorter100|6850_ , \new_Sorter100|6851_ ,
    \new_Sorter100|6852_ , \new_Sorter100|6853_ , \new_Sorter100|6854_ ,
    \new_Sorter100|6855_ , \new_Sorter100|6856_ , \new_Sorter100|6857_ ,
    \new_Sorter100|6858_ , \new_Sorter100|6859_ , \new_Sorter100|6860_ ,
    \new_Sorter100|6861_ , \new_Sorter100|6862_ , \new_Sorter100|6863_ ,
    \new_Sorter100|6864_ , \new_Sorter100|6865_ , \new_Sorter100|6866_ ,
    \new_Sorter100|6867_ , \new_Sorter100|6868_ , \new_Sorter100|6869_ ,
    \new_Sorter100|6870_ , \new_Sorter100|6871_ , \new_Sorter100|6872_ ,
    \new_Sorter100|6873_ , \new_Sorter100|6874_ , \new_Sorter100|6875_ ,
    \new_Sorter100|6876_ , \new_Sorter100|6877_ , \new_Sorter100|6878_ ,
    \new_Sorter100|6879_ , \new_Sorter100|6880_ , \new_Sorter100|6881_ ,
    \new_Sorter100|6882_ , \new_Sorter100|6883_ , \new_Sorter100|6884_ ,
    \new_Sorter100|6885_ , \new_Sorter100|6886_ , \new_Sorter100|6887_ ,
    \new_Sorter100|6888_ , \new_Sorter100|6889_ , \new_Sorter100|6890_ ,
    \new_Sorter100|6891_ , \new_Sorter100|6892_ , \new_Sorter100|6893_ ,
    \new_Sorter100|6894_ , \new_Sorter100|6895_ , \new_Sorter100|6896_ ,
    \new_Sorter100|6897_ , \new_Sorter100|6898_ , \new_Sorter100|6899_ ,
    \new_Sorter100|6900_ , \new_Sorter100|6999_ , \new_Sorter100|6901_ ,
    \new_Sorter100|6902_ , \new_Sorter100|6903_ , \new_Sorter100|6904_ ,
    \new_Sorter100|6905_ , \new_Sorter100|6906_ , \new_Sorter100|6907_ ,
    \new_Sorter100|6908_ , \new_Sorter100|6909_ , \new_Sorter100|6910_ ,
    \new_Sorter100|6911_ , \new_Sorter100|6912_ , \new_Sorter100|6913_ ,
    \new_Sorter100|6914_ , \new_Sorter100|6915_ , \new_Sorter100|6916_ ,
    \new_Sorter100|6917_ , \new_Sorter100|6918_ , \new_Sorter100|6919_ ,
    \new_Sorter100|6920_ , \new_Sorter100|6921_ , \new_Sorter100|6922_ ,
    \new_Sorter100|6923_ , \new_Sorter100|6924_ , \new_Sorter100|6925_ ,
    \new_Sorter100|6926_ , \new_Sorter100|6927_ , \new_Sorter100|6928_ ,
    \new_Sorter100|6929_ , \new_Sorter100|6930_ , \new_Sorter100|6931_ ,
    \new_Sorter100|6932_ , \new_Sorter100|6933_ , \new_Sorter100|6934_ ,
    \new_Sorter100|6935_ , \new_Sorter100|6936_ , \new_Sorter100|6937_ ,
    \new_Sorter100|6938_ , \new_Sorter100|6939_ , \new_Sorter100|6940_ ,
    \new_Sorter100|6941_ , \new_Sorter100|6942_ , \new_Sorter100|6943_ ,
    \new_Sorter100|6944_ , \new_Sorter100|6945_ , \new_Sorter100|6946_ ,
    \new_Sorter100|6947_ , \new_Sorter100|6948_ , \new_Sorter100|6949_ ,
    \new_Sorter100|6950_ , \new_Sorter100|6951_ , \new_Sorter100|6952_ ,
    \new_Sorter100|6953_ , \new_Sorter100|6954_ , \new_Sorter100|6955_ ,
    \new_Sorter100|6956_ , \new_Sorter100|6957_ , \new_Sorter100|6958_ ,
    \new_Sorter100|6959_ , \new_Sorter100|6960_ , \new_Sorter100|6961_ ,
    \new_Sorter100|6962_ , \new_Sorter100|6963_ , \new_Sorter100|6964_ ,
    \new_Sorter100|6965_ , \new_Sorter100|6966_ , \new_Sorter100|6967_ ,
    \new_Sorter100|6968_ , \new_Sorter100|6969_ , \new_Sorter100|6970_ ,
    \new_Sorter100|6971_ , \new_Sorter100|6972_ , \new_Sorter100|6973_ ,
    \new_Sorter100|6974_ , \new_Sorter100|6975_ , \new_Sorter100|6976_ ,
    \new_Sorter100|6977_ , \new_Sorter100|6978_ , \new_Sorter100|6979_ ,
    \new_Sorter100|6980_ , \new_Sorter100|6981_ , \new_Sorter100|6982_ ,
    \new_Sorter100|6983_ , \new_Sorter100|6984_ , \new_Sorter100|6985_ ,
    \new_Sorter100|6986_ , \new_Sorter100|6987_ , \new_Sorter100|6988_ ,
    \new_Sorter100|6989_ , \new_Sorter100|6990_ , \new_Sorter100|6991_ ,
    \new_Sorter100|6992_ , \new_Sorter100|6993_ , \new_Sorter100|6994_ ,
    \new_Sorter100|6995_ , \new_Sorter100|6996_ , \new_Sorter100|6997_ ,
    \new_Sorter100|6998_ , \new_Sorter100|7000_ , \new_Sorter100|7001_ ,
    \new_Sorter100|7002_ , \new_Sorter100|7003_ , \new_Sorter100|7004_ ,
    \new_Sorter100|7005_ , \new_Sorter100|7006_ , \new_Sorter100|7007_ ,
    \new_Sorter100|7008_ , \new_Sorter100|7009_ , \new_Sorter100|7010_ ,
    \new_Sorter100|7011_ , \new_Sorter100|7012_ , \new_Sorter100|7013_ ,
    \new_Sorter100|7014_ , \new_Sorter100|7015_ , \new_Sorter100|7016_ ,
    \new_Sorter100|7017_ , \new_Sorter100|7018_ , \new_Sorter100|7019_ ,
    \new_Sorter100|7020_ , \new_Sorter100|7021_ , \new_Sorter100|7022_ ,
    \new_Sorter100|7023_ , \new_Sorter100|7024_ , \new_Sorter100|7025_ ,
    \new_Sorter100|7026_ , \new_Sorter100|7027_ , \new_Sorter100|7028_ ,
    \new_Sorter100|7029_ , \new_Sorter100|7030_ , \new_Sorter100|7031_ ,
    \new_Sorter100|7032_ , \new_Sorter100|7033_ , \new_Sorter100|7034_ ,
    \new_Sorter100|7035_ , \new_Sorter100|7036_ , \new_Sorter100|7037_ ,
    \new_Sorter100|7038_ , \new_Sorter100|7039_ , \new_Sorter100|7040_ ,
    \new_Sorter100|7041_ , \new_Sorter100|7042_ , \new_Sorter100|7043_ ,
    \new_Sorter100|7044_ , \new_Sorter100|7045_ , \new_Sorter100|7046_ ,
    \new_Sorter100|7047_ , \new_Sorter100|7048_ , \new_Sorter100|7049_ ,
    \new_Sorter100|7050_ , \new_Sorter100|7051_ , \new_Sorter100|7052_ ,
    \new_Sorter100|7053_ , \new_Sorter100|7054_ , \new_Sorter100|7055_ ,
    \new_Sorter100|7056_ , \new_Sorter100|7057_ , \new_Sorter100|7058_ ,
    \new_Sorter100|7059_ , \new_Sorter100|7060_ , \new_Sorter100|7061_ ,
    \new_Sorter100|7062_ , \new_Sorter100|7063_ , \new_Sorter100|7064_ ,
    \new_Sorter100|7065_ , \new_Sorter100|7066_ , \new_Sorter100|7067_ ,
    \new_Sorter100|7068_ , \new_Sorter100|7069_ , \new_Sorter100|7070_ ,
    \new_Sorter100|7071_ , \new_Sorter100|7072_ , \new_Sorter100|7073_ ,
    \new_Sorter100|7074_ , \new_Sorter100|7075_ , \new_Sorter100|7076_ ,
    \new_Sorter100|7077_ , \new_Sorter100|7078_ , \new_Sorter100|7079_ ,
    \new_Sorter100|7080_ , \new_Sorter100|7081_ , \new_Sorter100|7082_ ,
    \new_Sorter100|7083_ , \new_Sorter100|7084_ , \new_Sorter100|7085_ ,
    \new_Sorter100|7086_ , \new_Sorter100|7087_ , \new_Sorter100|7088_ ,
    \new_Sorter100|7089_ , \new_Sorter100|7090_ , \new_Sorter100|7091_ ,
    \new_Sorter100|7092_ , \new_Sorter100|7093_ , \new_Sorter100|7094_ ,
    \new_Sorter100|7095_ , \new_Sorter100|7096_ , \new_Sorter100|7097_ ,
    \new_Sorter100|7098_ , \new_Sorter100|7099_ , \new_Sorter100|7100_ ,
    \new_Sorter100|7199_ , \new_Sorter100|7101_ , \new_Sorter100|7102_ ,
    \new_Sorter100|7103_ , \new_Sorter100|7104_ , \new_Sorter100|7105_ ,
    \new_Sorter100|7106_ , \new_Sorter100|7107_ , \new_Sorter100|7108_ ,
    \new_Sorter100|7109_ , \new_Sorter100|7110_ , \new_Sorter100|7111_ ,
    \new_Sorter100|7112_ , \new_Sorter100|7113_ , \new_Sorter100|7114_ ,
    \new_Sorter100|7115_ , \new_Sorter100|7116_ , \new_Sorter100|7117_ ,
    \new_Sorter100|7118_ , \new_Sorter100|7119_ , \new_Sorter100|7120_ ,
    \new_Sorter100|7121_ , \new_Sorter100|7122_ , \new_Sorter100|7123_ ,
    \new_Sorter100|7124_ , \new_Sorter100|7125_ , \new_Sorter100|7126_ ,
    \new_Sorter100|7127_ , \new_Sorter100|7128_ , \new_Sorter100|7129_ ,
    \new_Sorter100|7130_ , \new_Sorter100|7131_ , \new_Sorter100|7132_ ,
    \new_Sorter100|7133_ , \new_Sorter100|7134_ , \new_Sorter100|7135_ ,
    \new_Sorter100|7136_ , \new_Sorter100|7137_ , \new_Sorter100|7138_ ,
    \new_Sorter100|7139_ , \new_Sorter100|7140_ , \new_Sorter100|7141_ ,
    \new_Sorter100|7142_ , \new_Sorter100|7143_ , \new_Sorter100|7144_ ,
    \new_Sorter100|7145_ , \new_Sorter100|7146_ , \new_Sorter100|7147_ ,
    \new_Sorter100|7148_ , \new_Sorter100|7149_ , \new_Sorter100|7150_ ,
    \new_Sorter100|7151_ , \new_Sorter100|7152_ , \new_Sorter100|7153_ ,
    \new_Sorter100|7154_ , \new_Sorter100|7155_ , \new_Sorter100|7156_ ,
    \new_Sorter100|7157_ , \new_Sorter100|7158_ , \new_Sorter100|7159_ ,
    \new_Sorter100|7160_ , \new_Sorter100|7161_ , \new_Sorter100|7162_ ,
    \new_Sorter100|7163_ , \new_Sorter100|7164_ , \new_Sorter100|7165_ ,
    \new_Sorter100|7166_ , \new_Sorter100|7167_ , \new_Sorter100|7168_ ,
    \new_Sorter100|7169_ , \new_Sorter100|7170_ , \new_Sorter100|7171_ ,
    \new_Sorter100|7172_ , \new_Sorter100|7173_ , \new_Sorter100|7174_ ,
    \new_Sorter100|7175_ , \new_Sorter100|7176_ , \new_Sorter100|7177_ ,
    \new_Sorter100|7178_ , \new_Sorter100|7179_ , \new_Sorter100|7180_ ,
    \new_Sorter100|7181_ , \new_Sorter100|7182_ , \new_Sorter100|7183_ ,
    \new_Sorter100|7184_ , \new_Sorter100|7185_ , \new_Sorter100|7186_ ,
    \new_Sorter100|7187_ , \new_Sorter100|7188_ , \new_Sorter100|7189_ ,
    \new_Sorter100|7190_ , \new_Sorter100|7191_ , \new_Sorter100|7192_ ,
    \new_Sorter100|7193_ , \new_Sorter100|7194_ , \new_Sorter100|7195_ ,
    \new_Sorter100|7196_ , \new_Sorter100|7197_ , \new_Sorter100|7198_ ,
    \new_Sorter100|7200_ , \new_Sorter100|7201_ , \new_Sorter100|7202_ ,
    \new_Sorter100|7203_ , \new_Sorter100|7204_ , \new_Sorter100|7205_ ,
    \new_Sorter100|7206_ , \new_Sorter100|7207_ , \new_Sorter100|7208_ ,
    \new_Sorter100|7209_ , \new_Sorter100|7210_ , \new_Sorter100|7211_ ,
    \new_Sorter100|7212_ , \new_Sorter100|7213_ , \new_Sorter100|7214_ ,
    \new_Sorter100|7215_ , \new_Sorter100|7216_ , \new_Sorter100|7217_ ,
    \new_Sorter100|7218_ , \new_Sorter100|7219_ , \new_Sorter100|7220_ ,
    \new_Sorter100|7221_ , \new_Sorter100|7222_ , \new_Sorter100|7223_ ,
    \new_Sorter100|7224_ , \new_Sorter100|7225_ , \new_Sorter100|7226_ ,
    \new_Sorter100|7227_ , \new_Sorter100|7228_ , \new_Sorter100|7229_ ,
    \new_Sorter100|7230_ , \new_Sorter100|7231_ , \new_Sorter100|7232_ ,
    \new_Sorter100|7233_ , \new_Sorter100|7234_ , \new_Sorter100|7235_ ,
    \new_Sorter100|7236_ , \new_Sorter100|7237_ , \new_Sorter100|7238_ ,
    \new_Sorter100|7239_ , \new_Sorter100|7240_ , \new_Sorter100|7241_ ,
    \new_Sorter100|7242_ , \new_Sorter100|7243_ , \new_Sorter100|7244_ ,
    \new_Sorter100|7245_ , \new_Sorter100|7246_ , \new_Sorter100|7247_ ,
    \new_Sorter100|7248_ , \new_Sorter100|7249_ , \new_Sorter100|7250_ ,
    \new_Sorter100|7251_ , \new_Sorter100|7252_ , \new_Sorter100|7253_ ,
    \new_Sorter100|7254_ , \new_Sorter100|7255_ , \new_Sorter100|7256_ ,
    \new_Sorter100|7257_ , \new_Sorter100|7258_ , \new_Sorter100|7259_ ,
    \new_Sorter100|7260_ , \new_Sorter100|7261_ , \new_Sorter100|7262_ ,
    \new_Sorter100|7263_ , \new_Sorter100|7264_ , \new_Sorter100|7265_ ,
    \new_Sorter100|7266_ , \new_Sorter100|7267_ , \new_Sorter100|7268_ ,
    \new_Sorter100|7269_ , \new_Sorter100|7270_ , \new_Sorter100|7271_ ,
    \new_Sorter100|7272_ , \new_Sorter100|7273_ , \new_Sorter100|7274_ ,
    \new_Sorter100|7275_ , \new_Sorter100|7276_ , \new_Sorter100|7277_ ,
    \new_Sorter100|7278_ , \new_Sorter100|7279_ , \new_Sorter100|7280_ ,
    \new_Sorter100|7281_ , \new_Sorter100|7282_ , \new_Sorter100|7283_ ,
    \new_Sorter100|7284_ , \new_Sorter100|7285_ , \new_Sorter100|7286_ ,
    \new_Sorter100|7287_ , \new_Sorter100|7288_ , \new_Sorter100|7289_ ,
    \new_Sorter100|7290_ , \new_Sorter100|7291_ , \new_Sorter100|7292_ ,
    \new_Sorter100|7293_ , \new_Sorter100|7294_ , \new_Sorter100|7295_ ,
    \new_Sorter100|7296_ , \new_Sorter100|7297_ , \new_Sorter100|7298_ ,
    \new_Sorter100|7299_ , \new_Sorter100|7300_ , \new_Sorter100|7399_ ,
    \new_Sorter100|7301_ , \new_Sorter100|7302_ , \new_Sorter100|7303_ ,
    \new_Sorter100|7304_ , \new_Sorter100|7305_ , \new_Sorter100|7306_ ,
    \new_Sorter100|7307_ , \new_Sorter100|7308_ , \new_Sorter100|7309_ ,
    \new_Sorter100|7310_ , \new_Sorter100|7311_ , \new_Sorter100|7312_ ,
    \new_Sorter100|7313_ , \new_Sorter100|7314_ , \new_Sorter100|7315_ ,
    \new_Sorter100|7316_ , \new_Sorter100|7317_ , \new_Sorter100|7318_ ,
    \new_Sorter100|7319_ , \new_Sorter100|7320_ , \new_Sorter100|7321_ ,
    \new_Sorter100|7322_ , \new_Sorter100|7323_ , \new_Sorter100|7324_ ,
    \new_Sorter100|7325_ , \new_Sorter100|7326_ , \new_Sorter100|7327_ ,
    \new_Sorter100|7328_ , \new_Sorter100|7329_ , \new_Sorter100|7330_ ,
    \new_Sorter100|7331_ , \new_Sorter100|7332_ , \new_Sorter100|7333_ ,
    \new_Sorter100|7334_ , \new_Sorter100|7335_ , \new_Sorter100|7336_ ,
    \new_Sorter100|7337_ , \new_Sorter100|7338_ , \new_Sorter100|7339_ ,
    \new_Sorter100|7340_ , \new_Sorter100|7341_ , \new_Sorter100|7342_ ,
    \new_Sorter100|7343_ , \new_Sorter100|7344_ , \new_Sorter100|7345_ ,
    \new_Sorter100|7346_ , \new_Sorter100|7347_ , \new_Sorter100|7348_ ,
    \new_Sorter100|7349_ , \new_Sorter100|7350_ , \new_Sorter100|7351_ ,
    \new_Sorter100|7352_ , \new_Sorter100|7353_ , \new_Sorter100|7354_ ,
    \new_Sorter100|7355_ , \new_Sorter100|7356_ , \new_Sorter100|7357_ ,
    \new_Sorter100|7358_ , \new_Sorter100|7359_ , \new_Sorter100|7360_ ,
    \new_Sorter100|7361_ , \new_Sorter100|7362_ , \new_Sorter100|7363_ ,
    \new_Sorter100|7364_ , \new_Sorter100|7365_ , \new_Sorter100|7366_ ,
    \new_Sorter100|7367_ , \new_Sorter100|7368_ , \new_Sorter100|7369_ ,
    \new_Sorter100|7370_ , \new_Sorter100|7371_ , \new_Sorter100|7372_ ,
    \new_Sorter100|7373_ , \new_Sorter100|7374_ , \new_Sorter100|7375_ ,
    \new_Sorter100|7376_ , \new_Sorter100|7377_ , \new_Sorter100|7378_ ,
    \new_Sorter100|7379_ , \new_Sorter100|7380_ , \new_Sorter100|7381_ ,
    \new_Sorter100|7382_ , \new_Sorter100|7383_ , \new_Sorter100|7384_ ,
    \new_Sorter100|7385_ , \new_Sorter100|7386_ , \new_Sorter100|7387_ ,
    \new_Sorter100|7388_ , \new_Sorter100|7389_ , \new_Sorter100|7390_ ,
    \new_Sorter100|7391_ , \new_Sorter100|7392_ , \new_Sorter100|7393_ ,
    \new_Sorter100|7394_ , \new_Sorter100|7395_ , \new_Sorter100|7396_ ,
    \new_Sorter100|7397_ , \new_Sorter100|7398_ , \new_Sorter100|7400_ ,
    \new_Sorter100|7401_ , \new_Sorter100|7402_ , \new_Sorter100|7403_ ,
    \new_Sorter100|7404_ , \new_Sorter100|7405_ , \new_Sorter100|7406_ ,
    \new_Sorter100|7407_ , \new_Sorter100|7408_ , \new_Sorter100|7409_ ,
    \new_Sorter100|7410_ , \new_Sorter100|7411_ , \new_Sorter100|7412_ ,
    \new_Sorter100|7413_ , \new_Sorter100|7414_ , \new_Sorter100|7415_ ,
    \new_Sorter100|7416_ , \new_Sorter100|7417_ , \new_Sorter100|7418_ ,
    \new_Sorter100|7419_ , \new_Sorter100|7420_ , \new_Sorter100|7421_ ,
    \new_Sorter100|7422_ , \new_Sorter100|7423_ , \new_Sorter100|7424_ ,
    \new_Sorter100|7425_ , \new_Sorter100|7426_ , \new_Sorter100|7427_ ,
    \new_Sorter100|7428_ , \new_Sorter100|7429_ , \new_Sorter100|7430_ ,
    \new_Sorter100|7431_ , \new_Sorter100|7432_ , \new_Sorter100|7433_ ,
    \new_Sorter100|7434_ , \new_Sorter100|7435_ , \new_Sorter100|7436_ ,
    \new_Sorter100|7437_ , \new_Sorter100|7438_ , \new_Sorter100|7439_ ,
    \new_Sorter100|7440_ , \new_Sorter100|7441_ , \new_Sorter100|7442_ ,
    \new_Sorter100|7443_ , \new_Sorter100|7444_ , \new_Sorter100|7445_ ,
    \new_Sorter100|7446_ , \new_Sorter100|7447_ , \new_Sorter100|7448_ ,
    \new_Sorter100|7449_ , \new_Sorter100|7450_ , \new_Sorter100|7451_ ,
    \new_Sorter100|7452_ , \new_Sorter100|7453_ , \new_Sorter100|7454_ ,
    \new_Sorter100|7455_ , \new_Sorter100|7456_ , \new_Sorter100|7457_ ,
    \new_Sorter100|7458_ , \new_Sorter100|7459_ , \new_Sorter100|7460_ ,
    \new_Sorter100|7461_ , \new_Sorter100|7462_ , \new_Sorter100|7463_ ,
    \new_Sorter100|7464_ , \new_Sorter100|7465_ , \new_Sorter100|7466_ ,
    \new_Sorter100|7467_ , \new_Sorter100|7468_ , \new_Sorter100|7469_ ,
    \new_Sorter100|7470_ , \new_Sorter100|7471_ , \new_Sorter100|7472_ ,
    \new_Sorter100|7473_ , \new_Sorter100|7474_ , \new_Sorter100|7475_ ,
    \new_Sorter100|7476_ , \new_Sorter100|7477_ , \new_Sorter100|7478_ ,
    \new_Sorter100|7479_ , \new_Sorter100|7480_ , \new_Sorter100|7481_ ,
    \new_Sorter100|7482_ , \new_Sorter100|7483_ , \new_Sorter100|7484_ ,
    \new_Sorter100|7485_ , \new_Sorter100|7486_ , \new_Sorter100|7487_ ,
    \new_Sorter100|7488_ , \new_Sorter100|7489_ , \new_Sorter100|7490_ ,
    \new_Sorter100|7491_ , \new_Sorter100|7492_ , \new_Sorter100|7493_ ,
    \new_Sorter100|7494_ , \new_Sorter100|7495_ , \new_Sorter100|7496_ ,
    \new_Sorter100|7497_ , \new_Sorter100|7498_ , \new_Sorter100|7499_ ,
    \new_Sorter100|7500_ , \new_Sorter100|7599_ , \new_Sorter100|7501_ ,
    \new_Sorter100|7502_ , \new_Sorter100|7503_ , \new_Sorter100|7504_ ,
    \new_Sorter100|7505_ , \new_Sorter100|7506_ , \new_Sorter100|7507_ ,
    \new_Sorter100|7508_ , \new_Sorter100|7509_ , \new_Sorter100|7510_ ,
    \new_Sorter100|7511_ , \new_Sorter100|7512_ , \new_Sorter100|7513_ ,
    \new_Sorter100|7514_ , \new_Sorter100|7515_ , \new_Sorter100|7516_ ,
    \new_Sorter100|7517_ , \new_Sorter100|7518_ , \new_Sorter100|7519_ ,
    \new_Sorter100|7520_ , \new_Sorter100|7521_ , \new_Sorter100|7522_ ,
    \new_Sorter100|7523_ , \new_Sorter100|7524_ , \new_Sorter100|7525_ ,
    \new_Sorter100|7526_ , \new_Sorter100|7527_ , \new_Sorter100|7528_ ,
    \new_Sorter100|7529_ , \new_Sorter100|7530_ , \new_Sorter100|7531_ ,
    \new_Sorter100|7532_ , \new_Sorter100|7533_ , \new_Sorter100|7534_ ,
    \new_Sorter100|7535_ , \new_Sorter100|7536_ , \new_Sorter100|7537_ ,
    \new_Sorter100|7538_ , \new_Sorter100|7539_ , \new_Sorter100|7540_ ,
    \new_Sorter100|7541_ , \new_Sorter100|7542_ , \new_Sorter100|7543_ ,
    \new_Sorter100|7544_ , \new_Sorter100|7545_ , \new_Sorter100|7546_ ,
    \new_Sorter100|7547_ , \new_Sorter100|7548_ , \new_Sorter100|7549_ ,
    \new_Sorter100|7550_ , \new_Sorter100|7551_ , \new_Sorter100|7552_ ,
    \new_Sorter100|7553_ , \new_Sorter100|7554_ , \new_Sorter100|7555_ ,
    \new_Sorter100|7556_ , \new_Sorter100|7557_ , \new_Sorter100|7558_ ,
    \new_Sorter100|7559_ , \new_Sorter100|7560_ , \new_Sorter100|7561_ ,
    \new_Sorter100|7562_ , \new_Sorter100|7563_ , \new_Sorter100|7564_ ,
    \new_Sorter100|7565_ , \new_Sorter100|7566_ , \new_Sorter100|7567_ ,
    \new_Sorter100|7568_ , \new_Sorter100|7569_ , \new_Sorter100|7570_ ,
    \new_Sorter100|7571_ , \new_Sorter100|7572_ , \new_Sorter100|7573_ ,
    \new_Sorter100|7574_ , \new_Sorter100|7575_ , \new_Sorter100|7576_ ,
    \new_Sorter100|7577_ , \new_Sorter100|7578_ , \new_Sorter100|7579_ ,
    \new_Sorter100|7580_ , \new_Sorter100|7581_ , \new_Sorter100|7582_ ,
    \new_Sorter100|7583_ , \new_Sorter100|7584_ , \new_Sorter100|7585_ ,
    \new_Sorter100|7586_ , \new_Sorter100|7587_ , \new_Sorter100|7588_ ,
    \new_Sorter100|7589_ , \new_Sorter100|7590_ , \new_Sorter100|7591_ ,
    \new_Sorter100|7592_ , \new_Sorter100|7593_ , \new_Sorter100|7594_ ,
    \new_Sorter100|7595_ , \new_Sorter100|7596_ , \new_Sorter100|7597_ ,
    \new_Sorter100|7598_ , \new_Sorter100|7600_ , \new_Sorter100|7601_ ,
    \new_Sorter100|7602_ , \new_Sorter100|7603_ , \new_Sorter100|7604_ ,
    \new_Sorter100|7605_ , \new_Sorter100|7606_ , \new_Sorter100|7607_ ,
    \new_Sorter100|7608_ , \new_Sorter100|7609_ , \new_Sorter100|7610_ ,
    \new_Sorter100|7611_ , \new_Sorter100|7612_ , \new_Sorter100|7613_ ,
    \new_Sorter100|7614_ , \new_Sorter100|7615_ , \new_Sorter100|7616_ ,
    \new_Sorter100|7617_ , \new_Sorter100|7618_ , \new_Sorter100|7619_ ,
    \new_Sorter100|7620_ , \new_Sorter100|7621_ , \new_Sorter100|7622_ ,
    \new_Sorter100|7623_ , \new_Sorter100|7624_ , \new_Sorter100|7625_ ,
    \new_Sorter100|7626_ , \new_Sorter100|7627_ , \new_Sorter100|7628_ ,
    \new_Sorter100|7629_ , \new_Sorter100|7630_ , \new_Sorter100|7631_ ,
    \new_Sorter100|7632_ , \new_Sorter100|7633_ , \new_Sorter100|7634_ ,
    \new_Sorter100|7635_ , \new_Sorter100|7636_ , \new_Sorter100|7637_ ,
    \new_Sorter100|7638_ , \new_Sorter100|7639_ , \new_Sorter100|7640_ ,
    \new_Sorter100|7641_ , \new_Sorter100|7642_ , \new_Sorter100|7643_ ,
    \new_Sorter100|7644_ , \new_Sorter100|7645_ , \new_Sorter100|7646_ ,
    \new_Sorter100|7647_ , \new_Sorter100|7648_ , \new_Sorter100|7649_ ,
    \new_Sorter100|7650_ , \new_Sorter100|7651_ , \new_Sorter100|7652_ ,
    \new_Sorter100|7653_ , \new_Sorter100|7654_ , \new_Sorter100|7655_ ,
    \new_Sorter100|7656_ , \new_Sorter100|7657_ , \new_Sorter100|7658_ ,
    \new_Sorter100|7659_ , \new_Sorter100|7660_ , \new_Sorter100|7661_ ,
    \new_Sorter100|7662_ , \new_Sorter100|7663_ , \new_Sorter100|7664_ ,
    \new_Sorter100|7665_ , \new_Sorter100|7666_ , \new_Sorter100|7667_ ,
    \new_Sorter100|7668_ , \new_Sorter100|7669_ , \new_Sorter100|7670_ ,
    \new_Sorter100|7671_ , \new_Sorter100|7672_ , \new_Sorter100|7673_ ,
    \new_Sorter100|7674_ , \new_Sorter100|7675_ , \new_Sorter100|7676_ ,
    \new_Sorter100|7677_ , \new_Sorter100|7678_ , \new_Sorter100|7679_ ,
    \new_Sorter100|7680_ , \new_Sorter100|7681_ , \new_Sorter100|7682_ ,
    \new_Sorter100|7683_ , \new_Sorter100|7684_ , \new_Sorter100|7685_ ,
    \new_Sorter100|7686_ , \new_Sorter100|7687_ , \new_Sorter100|7688_ ,
    \new_Sorter100|7689_ , \new_Sorter100|7690_ , \new_Sorter100|7691_ ,
    \new_Sorter100|7692_ , \new_Sorter100|7693_ , \new_Sorter100|7694_ ,
    \new_Sorter100|7695_ , \new_Sorter100|7696_ , \new_Sorter100|7697_ ,
    \new_Sorter100|7698_ , \new_Sorter100|7699_ , \new_Sorter100|7700_ ,
    \new_Sorter100|7799_ , \new_Sorter100|7701_ , \new_Sorter100|7702_ ,
    \new_Sorter100|7703_ , \new_Sorter100|7704_ , \new_Sorter100|7705_ ,
    \new_Sorter100|7706_ , \new_Sorter100|7707_ , \new_Sorter100|7708_ ,
    \new_Sorter100|7709_ , \new_Sorter100|7710_ , \new_Sorter100|7711_ ,
    \new_Sorter100|7712_ , \new_Sorter100|7713_ , \new_Sorter100|7714_ ,
    \new_Sorter100|7715_ , \new_Sorter100|7716_ , \new_Sorter100|7717_ ,
    \new_Sorter100|7718_ , \new_Sorter100|7719_ , \new_Sorter100|7720_ ,
    \new_Sorter100|7721_ , \new_Sorter100|7722_ , \new_Sorter100|7723_ ,
    \new_Sorter100|7724_ , \new_Sorter100|7725_ , \new_Sorter100|7726_ ,
    \new_Sorter100|7727_ , \new_Sorter100|7728_ , \new_Sorter100|7729_ ,
    \new_Sorter100|7730_ , \new_Sorter100|7731_ , \new_Sorter100|7732_ ,
    \new_Sorter100|7733_ , \new_Sorter100|7734_ , \new_Sorter100|7735_ ,
    \new_Sorter100|7736_ , \new_Sorter100|7737_ , \new_Sorter100|7738_ ,
    \new_Sorter100|7739_ , \new_Sorter100|7740_ , \new_Sorter100|7741_ ,
    \new_Sorter100|7742_ , \new_Sorter100|7743_ , \new_Sorter100|7744_ ,
    \new_Sorter100|7745_ , \new_Sorter100|7746_ , \new_Sorter100|7747_ ,
    \new_Sorter100|7748_ , \new_Sorter100|7749_ , \new_Sorter100|7750_ ,
    \new_Sorter100|7751_ , \new_Sorter100|7752_ , \new_Sorter100|7753_ ,
    \new_Sorter100|7754_ , \new_Sorter100|7755_ , \new_Sorter100|7756_ ,
    \new_Sorter100|7757_ , \new_Sorter100|7758_ , \new_Sorter100|7759_ ,
    \new_Sorter100|7760_ , \new_Sorter100|7761_ , \new_Sorter100|7762_ ,
    \new_Sorter100|7763_ , \new_Sorter100|7764_ , \new_Sorter100|7765_ ,
    \new_Sorter100|7766_ , \new_Sorter100|7767_ , \new_Sorter100|7768_ ,
    \new_Sorter100|7769_ , \new_Sorter100|7770_ , \new_Sorter100|7771_ ,
    \new_Sorter100|7772_ , \new_Sorter100|7773_ , \new_Sorter100|7774_ ,
    \new_Sorter100|7775_ , \new_Sorter100|7776_ , \new_Sorter100|7777_ ,
    \new_Sorter100|7778_ , \new_Sorter100|7779_ , \new_Sorter100|7780_ ,
    \new_Sorter100|7781_ , \new_Sorter100|7782_ , \new_Sorter100|7783_ ,
    \new_Sorter100|7784_ , \new_Sorter100|7785_ , \new_Sorter100|7786_ ,
    \new_Sorter100|7787_ , \new_Sorter100|7788_ , \new_Sorter100|7789_ ,
    \new_Sorter100|7790_ , \new_Sorter100|7791_ , \new_Sorter100|7792_ ,
    \new_Sorter100|7793_ , \new_Sorter100|7794_ , \new_Sorter100|7795_ ,
    \new_Sorter100|7796_ , \new_Sorter100|7797_ , \new_Sorter100|7798_ ,
    \new_Sorter100|7800_ , \new_Sorter100|7801_ , \new_Sorter100|7802_ ,
    \new_Sorter100|7803_ , \new_Sorter100|7804_ , \new_Sorter100|7805_ ,
    \new_Sorter100|7806_ , \new_Sorter100|7807_ , \new_Sorter100|7808_ ,
    \new_Sorter100|7809_ , \new_Sorter100|7810_ , \new_Sorter100|7811_ ,
    \new_Sorter100|7812_ , \new_Sorter100|7813_ , \new_Sorter100|7814_ ,
    \new_Sorter100|7815_ , \new_Sorter100|7816_ , \new_Sorter100|7817_ ,
    \new_Sorter100|7818_ , \new_Sorter100|7819_ , \new_Sorter100|7820_ ,
    \new_Sorter100|7821_ , \new_Sorter100|7822_ , \new_Sorter100|7823_ ,
    \new_Sorter100|7824_ , \new_Sorter100|7825_ , \new_Sorter100|7826_ ,
    \new_Sorter100|7827_ , \new_Sorter100|7828_ , \new_Sorter100|7829_ ,
    \new_Sorter100|7830_ , \new_Sorter100|7831_ , \new_Sorter100|7832_ ,
    \new_Sorter100|7833_ , \new_Sorter100|7834_ , \new_Sorter100|7835_ ,
    \new_Sorter100|7836_ , \new_Sorter100|7837_ , \new_Sorter100|7838_ ,
    \new_Sorter100|7839_ , \new_Sorter100|7840_ , \new_Sorter100|7841_ ,
    \new_Sorter100|7842_ , \new_Sorter100|7843_ , \new_Sorter100|7844_ ,
    \new_Sorter100|7845_ , \new_Sorter100|7846_ , \new_Sorter100|7847_ ,
    \new_Sorter100|7848_ , \new_Sorter100|7849_ , \new_Sorter100|7850_ ,
    \new_Sorter100|7851_ , \new_Sorter100|7852_ , \new_Sorter100|7853_ ,
    \new_Sorter100|7854_ , \new_Sorter100|7855_ , \new_Sorter100|7856_ ,
    \new_Sorter100|7857_ , \new_Sorter100|7858_ , \new_Sorter100|7859_ ,
    \new_Sorter100|7860_ , \new_Sorter100|7861_ , \new_Sorter100|7862_ ,
    \new_Sorter100|7863_ , \new_Sorter100|7864_ , \new_Sorter100|7865_ ,
    \new_Sorter100|7866_ , \new_Sorter100|7867_ , \new_Sorter100|7868_ ,
    \new_Sorter100|7869_ , \new_Sorter100|7870_ , \new_Sorter100|7871_ ,
    \new_Sorter100|7872_ , \new_Sorter100|7873_ , \new_Sorter100|7874_ ,
    \new_Sorter100|7875_ , \new_Sorter100|7876_ , \new_Sorter100|7877_ ,
    \new_Sorter100|7878_ , \new_Sorter100|7879_ , \new_Sorter100|7880_ ,
    \new_Sorter100|7881_ , \new_Sorter100|7882_ , \new_Sorter100|7883_ ,
    \new_Sorter100|7884_ , \new_Sorter100|7885_ , \new_Sorter100|7886_ ,
    \new_Sorter100|7887_ , \new_Sorter100|7888_ , \new_Sorter100|7889_ ,
    \new_Sorter100|7890_ , \new_Sorter100|7891_ , \new_Sorter100|7892_ ,
    \new_Sorter100|7893_ , \new_Sorter100|7894_ , \new_Sorter100|7895_ ,
    \new_Sorter100|7896_ , \new_Sorter100|7897_ , \new_Sorter100|7898_ ,
    \new_Sorter100|7899_ , \new_Sorter100|7900_ , \new_Sorter100|7999_ ,
    \new_Sorter100|7901_ , \new_Sorter100|7902_ , \new_Sorter100|7903_ ,
    \new_Sorter100|7904_ , \new_Sorter100|7905_ , \new_Sorter100|7906_ ,
    \new_Sorter100|7907_ , \new_Sorter100|7908_ , \new_Sorter100|7909_ ,
    \new_Sorter100|7910_ , \new_Sorter100|7911_ , \new_Sorter100|7912_ ,
    \new_Sorter100|7913_ , \new_Sorter100|7914_ , \new_Sorter100|7915_ ,
    \new_Sorter100|7916_ , \new_Sorter100|7917_ , \new_Sorter100|7918_ ,
    \new_Sorter100|7919_ , \new_Sorter100|7920_ , \new_Sorter100|7921_ ,
    \new_Sorter100|7922_ , \new_Sorter100|7923_ , \new_Sorter100|7924_ ,
    \new_Sorter100|7925_ , \new_Sorter100|7926_ , \new_Sorter100|7927_ ,
    \new_Sorter100|7928_ , \new_Sorter100|7929_ , \new_Sorter100|7930_ ,
    \new_Sorter100|7931_ , \new_Sorter100|7932_ , \new_Sorter100|7933_ ,
    \new_Sorter100|7934_ , \new_Sorter100|7935_ , \new_Sorter100|7936_ ,
    \new_Sorter100|7937_ , \new_Sorter100|7938_ , \new_Sorter100|7939_ ,
    \new_Sorter100|7940_ , \new_Sorter100|7941_ , \new_Sorter100|7942_ ,
    \new_Sorter100|7943_ , \new_Sorter100|7944_ , \new_Sorter100|7945_ ,
    \new_Sorter100|7946_ , \new_Sorter100|7947_ , \new_Sorter100|7948_ ,
    \new_Sorter100|7949_ , \new_Sorter100|7950_ , \new_Sorter100|7951_ ,
    \new_Sorter100|7952_ , \new_Sorter100|7953_ , \new_Sorter100|7954_ ,
    \new_Sorter100|7955_ , \new_Sorter100|7956_ , \new_Sorter100|7957_ ,
    \new_Sorter100|7958_ , \new_Sorter100|7959_ , \new_Sorter100|7960_ ,
    \new_Sorter100|7961_ , \new_Sorter100|7962_ , \new_Sorter100|7963_ ,
    \new_Sorter100|7964_ , \new_Sorter100|7965_ , \new_Sorter100|7966_ ,
    \new_Sorter100|7967_ , \new_Sorter100|7968_ , \new_Sorter100|7969_ ,
    \new_Sorter100|7970_ , \new_Sorter100|7971_ , \new_Sorter100|7972_ ,
    \new_Sorter100|7973_ , \new_Sorter100|7974_ , \new_Sorter100|7975_ ,
    \new_Sorter100|7976_ , \new_Sorter100|7977_ , \new_Sorter100|7978_ ,
    \new_Sorter100|7979_ , \new_Sorter100|7980_ , \new_Sorter100|7981_ ,
    \new_Sorter100|7982_ , \new_Sorter100|7983_ , \new_Sorter100|7984_ ,
    \new_Sorter100|7985_ , \new_Sorter100|7986_ , \new_Sorter100|7987_ ,
    \new_Sorter100|7988_ , \new_Sorter100|7989_ , \new_Sorter100|7990_ ,
    \new_Sorter100|7991_ , \new_Sorter100|7992_ , \new_Sorter100|7993_ ,
    \new_Sorter100|7994_ , \new_Sorter100|7995_ , \new_Sorter100|7996_ ,
    \new_Sorter100|7997_ , \new_Sorter100|7998_ , \new_Sorter100|8000_ ,
    \new_Sorter100|8001_ , \new_Sorter100|8002_ , \new_Sorter100|8003_ ,
    \new_Sorter100|8004_ , \new_Sorter100|8005_ , \new_Sorter100|8006_ ,
    \new_Sorter100|8007_ , \new_Sorter100|8008_ , \new_Sorter100|8009_ ,
    \new_Sorter100|8010_ , \new_Sorter100|8011_ , \new_Sorter100|8012_ ,
    \new_Sorter100|8013_ , \new_Sorter100|8014_ , \new_Sorter100|8015_ ,
    \new_Sorter100|8016_ , \new_Sorter100|8017_ , \new_Sorter100|8018_ ,
    \new_Sorter100|8019_ , \new_Sorter100|8020_ , \new_Sorter100|8021_ ,
    \new_Sorter100|8022_ , \new_Sorter100|8023_ , \new_Sorter100|8024_ ,
    \new_Sorter100|8025_ , \new_Sorter100|8026_ , \new_Sorter100|8027_ ,
    \new_Sorter100|8028_ , \new_Sorter100|8029_ , \new_Sorter100|8030_ ,
    \new_Sorter100|8031_ , \new_Sorter100|8032_ , \new_Sorter100|8033_ ,
    \new_Sorter100|8034_ , \new_Sorter100|8035_ , \new_Sorter100|8036_ ,
    \new_Sorter100|8037_ , \new_Sorter100|8038_ , \new_Sorter100|8039_ ,
    \new_Sorter100|8040_ , \new_Sorter100|8041_ , \new_Sorter100|8042_ ,
    \new_Sorter100|8043_ , \new_Sorter100|8044_ , \new_Sorter100|8045_ ,
    \new_Sorter100|8046_ , \new_Sorter100|8047_ , \new_Sorter100|8048_ ,
    \new_Sorter100|8049_ , \new_Sorter100|8050_ , \new_Sorter100|8051_ ,
    \new_Sorter100|8052_ , \new_Sorter100|8053_ , \new_Sorter100|8054_ ,
    \new_Sorter100|8055_ , \new_Sorter100|8056_ , \new_Sorter100|8057_ ,
    \new_Sorter100|8058_ , \new_Sorter100|8059_ , \new_Sorter100|8060_ ,
    \new_Sorter100|8061_ , \new_Sorter100|8062_ , \new_Sorter100|8063_ ,
    \new_Sorter100|8064_ , \new_Sorter100|8065_ , \new_Sorter100|8066_ ,
    \new_Sorter100|8067_ , \new_Sorter100|8068_ , \new_Sorter100|8069_ ,
    \new_Sorter100|8070_ , \new_Sorter100|8071_ , \new_Sorter100|8072_ ,
    \new_Sorter100|8073_ , \new_Sorter100|8074_ , \new_Sorter100|8075_ ,
    \new_Sorter100|8076_ , \new_Sorter100|8077_ , \new_Sorter100|8078_ ,
    \new_Sorter100|8079_ , \new_Sorter100|8080_ , \new_Sorter100|8081_ ,
    \new_Sorter100|8082_ , \new_Sorter100|8083_ , \new_Sorter100|8084_ ,
    \new_Sorter100|8085_ , \new_Sorter100|8086_ , \new_Sorter100|8087_ ,
    \new_Sorter100|8088_ , \new_Sorter100|8089_ , \new_Sorter100|8090_ ,
    \new_Sorter100|8091_ , \new_Sorter100|8092_ , \new_Sorter100|8093_ ,
    \new_Sorter100|8094_ , \new_Sorter100|8095_ , \new_Sorter100|8096_ ,
    \new_Sorter100|8097_ , \new_Sorter100|8098_ , \new_Sorter100|8099_ ,
    \new_Sorter100|8100_ , \new_Sorter100|8199_ , \new_Sorter100|8101_ ,
    \new_Sorter100|8102_ , \new_Sorter100|8103_ , \new_Sorter100|8104_ ,
    \new_Sorter100|8105_ , \new_Sorter100|8106_ , \new_Sorter100|8107_ ,
    \new_Sorter100|8108_ , \new_Sorter100|8109_ , \new_Sorter100|8110_ ,
    \new_Sorter100|8111_ , \new_Sorter100|8112_ , \new_Sorter100|8113_ ,
    \new_Sorter100|8114_ , \new_Sorter100|8115_ , \new_Sorter100|8116_ ,
    \new_Sorter100|8117_ , \new_Sorter100|8118_ , \new_Sorter100|8119_ ,
    \new_Sorter100|8120_ , \new_Sorter100|8121_ , \new_Sorter100|8122_ ,
    \new_Sorter100|8123_ , \new_Sorter100|8124_ , \new_Sorter100|8125_ ,
    \new_Sorter100|8126_ , \new_Sorter100|8127_ , \new_Sorter100|8128_ ,
    \new_Sorter100|8129_ , \new_Sorter100|8130_ , \new_Sorter100|8131_ ,
    \new_Sorter100|8132_ , \new_Sorter100|8133_ , \new_Sorter100|8134_ ,
    \new_Sorter100|8135_ , \new_Sorter100|8136_ , \new_Sorter100|8137_ ,
    \new_Sorter100|8138_ , \new_Sorter100|8139_ , \new_Sorter100|8140_ ,
    \new_Sorter100|8141_ , \new_Sorter100|8142_ , \new_Sorter100|8143_ ,
    \new_Sorter100|8144_ , \new_Sorter100|8145_ , \new_Sorter100|8146_ ,
    \new_Sorter100|8147_ , \new_Sorter100|8148_ , \new_Sorter100|8149_ ,
    \new_Sorter100|8150_ , \new_Sorter100|8151_ , \new_Sorter100|8152_ ,
    \new_Sorter100|8153_ , \new_Sorter100|8154_ , \new_Sorter100|8155_ ,
    \new_Sorter100|8156_ , \new_Sorter100|8157_ , \new_Sorter100|8158_ ,
    \new_Sorter100|8159_ , \new_Sorter100|8160_ , \new_Sorter100|8161_ ,
    \new_Sorter100|8162_ , \new_Sorter100|8163_ , \new_Sorter100|8164_ ,
    \new_Sorter100|8165_ , \new_Sorter100|8166_ , \new_Sorter100|8167_ ,
    \new_Sorter100|8168_ , \new_Sorter100|8169_ , \new_Sorter100|8170_ ,
    \new_Sorter100|8171_ , \new_Sorter100|8172_ , \new_Sorter100|8173_ ,
    \new_Sorter100|8174_ , \new_Sorter100|8175_ , \new_Sorter100|8176_ ,
    \new_Sorter100|8177_ , \new_Sorter100|8178_ , \new_Sorter100|8179_ ,
    \new_Sorter100|8180_ , \new_Sorter100|8181_ , \new_Sorter100|8182_ ,
    \new_Sorter100|8183_ , \new_Sorter100|8184_ , \new_Sorter100|8185_ ,
    \new_Sorter100|8186_ , \new_Sorter100|8187_ , \new_Sorter100|8188_ ,
    \new_Sorter100|8189_ , \new_Sorter100|8190_ , \new_Sorter100|8191_ ,
    \new_Sorter100|8192_ , \new_Sorter100|8193_ , \new_Sorter100|8194_ ,
    \new_Sorter100|8195_ , \new_Sorter100|8196_ , \new_Sorter100|8197_ ,
    \new_Sorter100|8198_ , \new_Sorter100|8200_ , \new_Sorter100|8201_ ,
    \new_Sorter100|8202_ , \new_Sorter100|8203_ , \new_Sorter100|8204_ ,
    \new_Sorter100|8205_ , \new_Sorter100|8206_ , \new_Sorter100|8207_ ,
    \new_Sorter100|8208_ , \new_Sorter100|8209_ , \new_Sorter100|8210_ ,
    \new_Sorter100|8211_ , \new_Sorter100|8212_ , \new_Sorter100|8213_ ,
    \new_Sorter100|8214_ , \new_Sorter100|8215_ , \new_Sorter100|8216_ ,
    \new_Sorter100|8217_ , \new_Sorter100|8218_ , \new_Sorter100|8219_ ,
    \new_Sorter100|8220_ , \new_Sorter100|8221_ , \new_Sorter100|8222_ ,
    \new_Sorter100|8223_ , \new_Sorter100|8224_ , \new_Sorter100|8225_ ,
    \new_Sorter100|8226_ , \new_Sorter100|8227_ , \new_Sorter100|8228_ ,
    \new_Sorter100|8229_ , \new_Sorter100|8230_ , \new_Sorter100|8231_ ,
    \new_Sorter100|8232_ , \new_Sorter100|8233_ , \new_Sorter100|8234_ ,
    \new_Sorter100|8235_ , \new_Sorter100|8236_ , \new_Sorter100|8237_ ,
    \new_Sorter100|8238_ , \new_Sorter100|8239_ , \new_Sorter100|8240_ ,
    \new_Sorter100|8241_ , \new_Sorter100|8242_ , \new_Sorter100|8243_ ,
    \new_Sorter100|8244_ , \new_Sorter100|8245_ , \new_Sorter100|8246_ ,
    \new_Sorter100|8247_ , \new_Sorter100|8248_ , \new_Sorter100|8249_ ,
    \new_Sorter100|8250_ , \new_Sorter100|8251_ , \new_Sorter100|8252_ ,
    \new_Sorter100|8253_ , \new_Sorter100|8254_ , \new_Sorter100|8255_ ,
    \new_Sorter100|8256_ , \new_Sorter100|8257_ , \new_Sorter100|8258_ ,
    \new_Sorter100|8259_ , \new_Sorter100|8260_ , \new_Sorter100|8261_ ,
    \new_Sorter100|8262_ , \new_Sorter100|8263_ , \new_Sorter100|8264_ ,
    \new_Sorter100|8265_ , \new_Sorter100|8266_ , \new_Sorter100|8267_ ,
    \new_Sorter100|8268_ , \new_Sorter100|8269_ , \new_Sorter100|8270_ ,
    \new_Sorter100|8271_ , \new_Sorter100|8272_ , \new_Sorter100|8273_ ,
    \new_Sorter100|8274_ , \new_Sorter100|8275_ , \new_Sorter100|8276_ ,
    \new_Sorter100|8277_ , \new_Sorter100|8278_ , \new_Sorter100|8279_ ,
    \new_Sorter100|8280_ , \new_Sorter100|8281_ , \new_Sorter100|8282_ ,
    \new_Sorter100|8283_ , \new_Sorter100|8284_ , \new_Sorter100|8285_ ,
    \new_Sorter100|8286_ , \new_Sorter100|8287_ , \new_Sorter100|8288_ ,
    \new_Sorter100|8289_ , \new_Sorter100|8290_ , \new_Sorter100|8291_ ,
    \new_Sorter100|8292_ , \new_Sorter100|8293_ , \new_Sorter100|8294_ ,
    \new_Sorter100|8295_ , \new_Sorter100|8296_ , \new_Sorter100|8297_ ,
    \new_Sorter100|8298_ , \new_Sorter100|8299_ , \new_Sorter100|8300_ ,
    \new_Sorter100|8399_ , \new_Sorter100|8301_ , \new_Sorter100|8302_ ,
    \new_Sorter100|8303_ , \new_Sorter100|8304_ , \new_Sorter100|8305_ ,
    \new_Sorter100|8306_ , \new_Sorter100|8307_ , \new_Sorter100|8308_ ,
    \new_Sorter100|8309_ , \new_Sorter100|8310_ , \new_Sorter100|8311_ ,
    \new_Sorter100|8312_ , \new_Sorter100|8313_ , \new_Sorter100|8314_ ,
    \new_Sorter100|8315_ , \new_Sorter100|8316_ , \new_Sorter100|8317_ ,
    \new_Sorter100|8318_ , \new_Sorter100|8319_ , \new_Sorter100|8320_ ,
    \new_Sorter100|8321_ , \new_Sorter100|8322_ , \new_Sorter100|8323_ ,
    \new_Sorter100|8324_ , \new_Sorter100|8325_ , \new_Sorter100|8326_ ,
    \new_Sorter100|8327_ , \new_Sorter100|8328_ , \new_Sorter100|8329_ ,
    \new_Sorter100|8330_ , \new_Sorter100|8331_ , \new_Sorter100|8332_ ,
    \new_Sorter100|8333_ , \new_Sorter100|8334_ , \new_Sorter100|8335_ ,
    \new_Sorter100|8336_ , \new_Sorter100|8337_ , \new_Sorter100|8338_ ,
    \new_Sorter100|8339_ , \new_Sorter100|8340_ , \new_Sorter100|8341_ ,
    \new_Sorter100|8342_ , \new_Sorter100|8343_ , \new_Sorter100|8344_ ,
    \new_Sorter100|8345_ , \new_Sorter100|8346_ , \new_Sorter100|8347_ ,
    \new_Sorter100|8348_ , \new_Sorter100|8349_ , \new_Sorter100|8350_ ,
    \new_Sorter100|8351_ , \new_Sorter100|8352_ , \new_Sorter100|8353_ ,
    \new_Sorter100|8354_ , \new_Sorter100|8355_ , \new_Sorter100|8356_ ,
    \new_Sorter100|8357_ , \new_Sorter100|8358_ , \new_Sorter100|8359_ ,
    \new_Sorter100|8360_ , \new_Sorter100|8361_ , \new_Sorter100|8362_ ,
    \new_Sorter100|8363_ , \new_Sorter100|8364_ , \new_Sorter100|8365_ ,
    \new_Sorter100|8366_ , \new_Sorter100|8367_ , \new_Sorter100|8368_ ,
    \new_Sorter100|8369_ , \new_Sorter100|8370_ , \new_Sorter100|8371_ ,
    \new_Sorter100|8372_ , \new_Sorter100|8373_ , \new_Sorter100|8374_ ,
    \new_Sorter100|8375_ , \new_Sorter100|8376_ , \new_Sorter100|8377_ ,
    \new_Sorter100|8378_ , \new_Sorter100|8379_ , \new_Sorter100|8380_ ,
    \new_Sorter100|8381_ , \new_Sorter100|8382_ , \new_Sorter100|8383_ ,
    \new_Sorter100|8384_ , \new_Sorter100|8385_ , \new_Sorter100|8386_ ,
    \new_Sorter100|8387_ , \new_Sorter100|8388_ , \new_Sorter100|8389_ ,
    \new_Sorter100|8390_ , \new_Sorter100|8391_ , \new_Sorter100|8392_ ,
    \new_Sorter100|8393_ , \new_Sorter100|8394_ , \new_Sorter100|8395_ ,
    \new_Sorter100|8396_ , \new_Sorter100|8397_ , \new_Sorter100|8398_ ,
    \new_Sorter100|8400_ , \new_Sorter100|8401_ , \new_Sorter100|8402_ ,
    \new_Sorter100|8403_ , \new_Sorter100|8404_ , \new_Sorter100|8405_ ,
    \new_Sorter100|8406_ , \new_Sorter100|8407_ , \new_Sorter100|8408_ ,
    \new_Sorter100|8409_ , \new_Sorter100|8410_ , \new_Sorter100|8411_ ,
    \new_Sorter100|8412_ , \new_Sorter100|8413_ , \new_Sorter100|8414_ ,
    \new_Sorter100|8415_ , \new_Sorter100|8416_ , \new_Sorter100|8417_ ,
    \new_Sorter100|8418_ , \new_Sorter100|8419_ , \new_Sorter100|8420_ ,
    \new_Sorter100|8421_ , \new_Sorter100|8422_ , \new_Sorter100|8423_ ,
    \new_Sorter100|8424_ , \new_Sorter100|8425_ , \new_Sorter100|8426_ ,
    \new_Sorter100|8427_ , \new_Sorter100|8428_ , \new_Sorter100|8429_ ,
    \new_Sorter100|8430_ , \new_Sorter100|8431_ , \new_Sorter100|8432_ ,
    \new_Sorter100|8433_ , \new_Sorter100|8434_ , \new_Sorter100|8435_ ,
    \new_Sorter100|8436_ , \new_Sorter100|8437_ , \new_Sorter100|8438_ ,
    \new_Sorter100|8439_ , \new_Sorter100|8440_ , \new_Sorter100|8441_ ,
    \new_Sorter100|8442_ , \new_Sorter100|8443_ , \new_Sorter100|8444_ ,
    \new_Sorter100|8445_ , \new_Sorter100|8446_ , \new_Sorter100|8447_ ,
    \new_Sorter100|8448_ , \new_Sorter100|8449_ , \new_Sorter100|8450_ ,
    \new_Sorter100|8451_ , \new_Sorter100|8452_ , \new_Sorter100|8453_ ,
    \new_Sorter100|8454_ , \new_Sorter100|8455_ , \new_Sorter100|8456_ ,
    \new_Sorter100|8457_ , \new_Sorter100|8458_ , \new_Sorter100|8459_ ,
    \new_Sorter100|8460_ , \new_Sorter100|8461_ , \new_Sorter100|8462_ ,
    \new_Sorter100|8463_ , \new_Sorter100|8464_ , \new_Sorter100|8465_ ,
    \new_Sorter100|8466_ , \new_Sorter100|8467_ , \new_Sorter100|8468_ ,
    \new_Sorter100|8469_ , \new_Sorter100|8470_ , \new_Sorter100|8471_ ,
    \new_Sorter100|8472_ , \new_Sorter100|8473_ , \new_Sorter100|8474_ ,
    \new_Sorter100|8475_ , \new_Sorter100|8476_ , \new_Sorter100|8477_ ,
    \new_Sorter100|8478_ , \new_Sorter100|8479_ , \new_Sorter100|8480_ ,
    \new_Sorter100|8481_ , \new_Sorter100|8482_ , \new_Sorter100|8483_ ,
    \new_Sorter100|8484_ , \new_Sorter100|8485_ , \new_Sorter100|8486_ ,
    \new_Sorter100|8487_ , \new_Sorter100|8488_ , \new_Sorter100|8489_ ,
    \new_Sorter100|8490_ , \new_Sorter100|8491_ , \new_Sorter100|8492_ ,
    \new_Sorter100|8493_ , \new_Sorter100|8494_ , \new_Sorter100|8495_ ,
    \new_Sorter100|8496_ , \new_Sorter100|8497_ , \new_Sorter100|8498_ ,
    \new_Sorter100|8499_ , \new_Sorter100|8500_ , \new_Sorter100|8599_ ,
    \new_Sorter100|8501_ , \new_Sorter100|8502_ , \new_Sorter100|8503_ ,
    \new_Sorter100|8504_ , \new_Sorter100|8505_ , \new_Sorter100|8506_ ,
    \new_Sorter100|8507_ , \new_Sorter100|8508_ , \new_Sorter100|8509_ ,
    \new_Sorter100|8510_ , \new_Sorter100|8511_ , \new_Sorter100|8512_ ,
    \new_Sorter100|8513_ , \new_Sorter100|8514_ , \new_Sorter100|8515_ ,
    \new_Sorter100|8516_ , \new_Sorter100|8517_ , \new_Sorter100|8518_ ,
    \new_Sorter100|8519_ , \new_Sorter100|8520_ , \new_Sorter100|8521_ ,
    \new_Sorter100|8522_ , \new_Sorter100|8523_ , \new_Sorter100|8524_ ,
    \new_Sorter100|8525_ , \new_Sorter100|8526_ , \new_Sorter100|8527_ ,
    \new_Sorter100|8528_ , \new_Sorter100|8529_ , \new_Sorter100|8530_ ,
    \new_Sorter100|8531_ , \new_Sorter100|8532_ , \new_Sorter100|8533_ ,
    \new_Sorter100|8534_ , \new_Sorter100|8535_ , \new_Sorter100|8536_ ,
    \new_Sorter100|8537_ , \new_Sorter100|8538_ , \new_Sorter100|8539_ ,
    \new_Sorter100|8540_ , \new_Sorter100|8541_ , \new_Sorter100|8542_ ,
    \new_Sorter100|8543_ , \new_Sorter100|8544_ , \new_Sorter100|8545_ ,
    \new_Sorter100|8546_ , \new_Sorter100|8547_ , \new_Sorter100|8548_ ,
    \new_Sorter100|8549_ , \new_Sorter100|8550_ , \new_Sorter100|8551_ ,
    \new_Sorter100|8552_ , \new_Sorter100|8553_ , \new_Sorter100|8554_ ,
    \new_Sorter100|8555_ , \new_Sorter100|8556_ , \new_Sorter100|8557_ ,
    \new_Sorter100|8558_ , \new_Sorter100|8559_ , \new_Sorter100|8560_ ,
    \new_Sorter100|8561_ , \new_Sorter100|8562_ , \new_Sorter100|8563_ ,
    \new_Sorter100|8564_ , \new_Sorter100|8565_ , \new_Sorter100|8566_ ,
    \new_Sorter100|8567_ , \new_Sorter100|8568_ , \new_Sorter100|8569_ ,
    \new_Sorter100|8570_ , \new_Sorter100|8571_ , \new_Sorter100|8572_ ,
    \new_Sorter100|8573_ , \new_Sorter100|8574_ , \new_Sorter100|8575_ ,
    \new_Sorter100|8576_ , \new_Sorter100|8577_ , \new_Sorter100|8578_ ,
    \new_Sorter100|8579_ , \new_Sorter100|8580_ , \new_Sorter100|8581_ ,
    \new_Sorter100|8582_ , \new_Sorter100|8583_ , \new_Sorter100|8584_ ,
    \new_Sorter100|8585_ , \new_Sorter100|8586_ , \new_Sorter100|8587_ ,
    \new_Sorter100|8588_ , \new_Sorter100|8589_ , \new_Sorter100|8590_ ,
    \new_Sorter100|8591_ , \new_Sorter100|8592_ , \new_Sorter100|8593_ ,
    \new_Sorter100|8594_ , \new_Sorter100|8595_ , \new_Sorter100|8596_ ,
    \new_Sorter100|8597_ , \new_Sorter100|8598_ , \new_Sorter100|8600_ ,
    \new_Sorter100|8601_ , \new_Sorter100|8602_ , \new_Sorter100|8603_ ,
    \new_Sorter100|8604_ , \new_Sorter100|8605_ , \new_Sorter100|8606_ ,
    \new_Sorter100|8607_ , \new_Sorter100|8608_ , \new_Sorter100|8609_ ,
    \new_Sorter100|8610_ , \new_Sorter100|8611_ , \new_Sorter100|8612_ ,
    \new_Sorter100|8613_ , \new_Sorter100|8614_ , \new_Sorter100|8615_ ,
    \new_Sorter100|8616_ , \new_Sorter100|8617_ , \new_Sorter100|8618_ ,
    \new_Sorter100|8619_ , \new_Sorter100|8620_ , \new_Sorter100|8621_ ,
    \new_Sorter100|8622_ , \new_Sorter100|8623_ , \new_Sorter100|8624_ ,
    \new_Sorter100|8625_ , \new_Sorter100|8626_ , \new_Sorter100|8627_ ,
    \new_Sorter100|8628_ , \new_Sorter100|8629_ , \new_Sorter100|8630_ ,
    \new_Sorter100|8631_ , \new_Sorter100|8632_ , \new_Sorter100|8633_ ,
    \new_Sorter100|8634_ , \new_Sorter100|8635_ , \new_Sorter100|8636_ ,
    \new_Sorter100|8637_ , \new_Sorter100|8638_ , \new_Sorter100|8639_ ,
    \new_Sorter100|8640_ , \new_Sorter100|8641_ , \new_Sorter100|8642_ ,
    \new_Sorter100|8643_ , \new_Sorter100|8644_ , \new_Sorter100|8645_ ,
    \new_Sorter100|8646_ , \new_Sorter100|8647_ , \new_Sorter100|8648_ ,
    \new_Sorter100|8649_ , \new_Sorter100|8650_ , \new_Sorter100|8651_ ,
    \new_Sorter100|8652_ , \new_Sorter100|8653_ , \new_Sorter100|8654_ ,
    \new_Sorter100|8655_ , \new_Sorter100|8656_ , \new_Sorter100|8657_ ,
    \new_Sorter100|8658_ , \new_Sorter100|8659_ , \new_Sorter100|8660_ ,
    \new_Sorter100|8661_ , \new_Sorter100|8662_ , \new_Sorter100|8663_ ,
    \new_Sorter100|8664_ , \new_Sorter100|8665_ , \new_Sorter100|8666_ ,
    \new_Sorter100|8667_ , \new_Sorter100|8668_ , \new_Sorter100|8669_ ,
    \new_Sorter100|8670_ , \new_Sorter100|8671_ , \new_Sorter100|8672_ ,
    \new_Sorter100|8673_ , \new_Sorter100|8674_ , \new_Sorter100|8675_ ,
    \new_Sorter100|8676_ , \new_Sorter100|8677_ , \new_Sorter100|8678_ ,
    \new_Sorter100|8679_ , \new_Sorter100|8680_ , \new_Sorter100|8681_ ,
    \new_Sorter100|8682_ , \new_Sorter100|8683_ , \new_Sorter100|8684_ ,
    \new_Sorter100|8685_ , \new_Sorter100|8686_ , \new_Sorter100|8687_ ,
    \new_Sorter100|8688_ , \new_Sorter100|8689_ , \new_Sorter100|8690_ ,
    \new_Sorter100|8691_ , \new_Sorter100|8692_ , \new_Sorter100|8693_ ,
    \new_Sorter100|8694_ , \new_Sorter100|8695_ , \new_Sorter100|8696_ ,
    \new_Sorter100|8697_ , \new_Sorter100|8698_ , \new_Sorter100|8699_ ,
    \new_Sorter100|8700_ , \new_Sorter100|8799_ , \new_Sorter100|8701_ ,
    \new_Sorter100|8702_ , \new_Sorter100|8703_ , \new_Sorter100|8704_ ,
    \new_Sorter100|8705_ , \new_Sorter100|8706_ , \new_Sorter100|8707_ ,
    \new_Sorter100|8708_ , \new_Sorter100|8709_ , \new_Sorter100|8710_ ,
    \new_Sorter100|8711_ , \new_Sorter100|8712_ , \new_Sorter100|8713_ ,
    \new_Sorter100|8714_ , \new_Sorter100|8715_ , \new_Sorter100|8716_ ,
    \new_Sorter100|8717_ , \new_Sorter100|8718_ , \new_Sorter100|8719_ ,
    \new_Sorter100|8720_ , \new_Sorter100|8721_ , \new_Sorter100|8722_ ,
    \new_Sorter100|8723_ , \new_Sorter100|8724_ , \new_Sorter100|8725_ ,
    \new_Sorter100|8726_ , \new_Sorter100|8727_ , \new_Sorter100|8728_ ,
    \new_Sorter100|8729_ , \new_Sorter100|8730_ , \new_Sorter100|8731_ ,
    \new_Sorter100|8732_ , \new_Sorter100|8733_ , \new_Sorter100|8734_ ,
    \new_Sorter100|8735_ , \new_Sorter100|8736_ , \new_Sorter100|8737_ ,
    \new_Sorter100|8738_ , \new_Sorter100|8739_ , \new_Sorter100|8740_ ,
    \new_Sorter100|8741_ , \new_Sorter100|8742_ , \new_Sorter100|8743_ ,
    \new_Sorter100|8744_ , \new_Sorter100|8745_ , \new_Sorter100|8746_ ,
    \new_Sorter100|8747_ , \new_Sorter100|8748_ , \new_Sorter100|8749_ ,
    \new_Sorter100|8750_ , \new_Sorter100|8751_ , \new_Sorter100|8752_ ,
    \new_Sorter100|8753_ , \new_Sorter100|8754_ , \new_Sorter100|8755_ ,
    \new_Sorter100|8756_ , \new_Sorter100|8757_ , \new_Sorter100|8758_ ,
    \new_Sorter100|8759_ , \new_Sorter100|8760_ , \new_Sorter100|8761_ ,
    \new_Sorter100|8762_ , \new_Sorter100|8763_ , \new_Sorter100|8764_ ,
    \new_Sorter100|8765_ , \new_Sorter100|8766_ , \new_Sorter100|8767_ ,
    \new_Sorter100|8768_ , \new_Sorter100|8769_ , \new_Sorter100|8770_ ,
    \new_Sorter100|8771_ , \new_Sorter100|8772_ , \new_Sorter100|8773_ ,
    \new_Sorter100|8774_ , \new_Sorter100|8775_ , \new_Sorter100|8776_ ,
    \new_Sorter100|8777_ , \new_Sorter100|8778_ , \new_Sorter100|8779_ ,
    \new_Sorter100|8780_ , \new_Sorter100|8781_ , \new_Sorter100|8782_ ,
    \new_Sorter100|8783_ , \new_Sorter100|8784_ , \new_Sorter100|8785_ ,
    \new_Sorter100|8786_ , \new_Sorter100|8787_ , \new_Sorter100|8788_ ,
    \new_Sorter100|8789_ , \new_Sorter100|8790_ , \new_Sorter100|8791_ ,
    \new_Sorter100|8792_ , \new_Sorter100|8793_ , \new_Sorter100|8794_ ,
    \new_Sorter100|8795_ , \new_Sorter100|8796_ , \new_Sorter100|8797_ ,
    \new_Sorter100|8798_ , \new_Sorter100|8800_ , \new_Sorter100|8801_ ,
    \new_Sorter100|8802_ , \new_Sorter100|8803_ , \new_Sorter100|8804_ ,
    \new_Sorter100|8805_ , \new_Sorter100|8806_ , \new_Sorter100|8807_ ,
    \new_Sorter100|8808_ , \new_Sorter100|8809_ , \new_Sorter100|8810_ ,
    \new_Sorter100|8811_ , \new_Sorter100|8812_ , \new_Sorter100|8813_ ,
    \new_Sorter100|8814_ , \new_Sorter100|8815_ , \new_Sorter100|8816_ ,
    \new_Sorter100|8817_ , \new_Sorter100|8818_ , \new_Sorter100|8819_ ,
    \new_Sorter100|8820_ , \new_Sorter100|8821_ , \new_Sorter100|8822_ ,
    \new_Sorter100|8823_ , \new_Sorter100|8824_ , \new_Sorter100|8825_ ,
    \new_Sorter100|8826_ , \new_Sorter100|8827_ , \new_Sorter100|8828_ ,
    \new_Sorter100|8829_ , \new_Sorter100|8830_ , \new_Sorter100|8831_ ,
    \new_Sorter100|8832_ , \new_Sorter100|8833_ , \new_Sorter100|8834_ ,
    \new_Sorter100|8835_ , \new_Sorter100|8836_ , \new_Sorter100|8837_ ,
    \new_Sorter100|8838_ , \new_Sorter100|8839_ , \new_Sorter100|8840_ ,
    \new_Sorter100|8841_ , \new_Sorter100|8842_ , \new_Sorter100|8843_ ,
    \new_Sorter100|8844_ , \new_Sorter100|8845_ , \new_Sorter100|8846_ ,
    \new_Sorter100|8847_ , \new_Sorter100|8848_ , \new_Sorter100|8849_ ,
    \new_Sorter100|8850_ , \new_Sorter100|8851_ , \new_Sorter100|8852_ ,
    \new_Sorter100|8853_ , \new_Sorter100|8854_ , \new_Sorter100|8855_ ,
    \new_Sorter100|8856_ , \new_Sorter100|8857_ , \new_Sorter100|8858_ ,
    \new_Sorter100|8859_ , \new_Sorter100|8860_ , \new_Sorter100|8861_ ,
    \new_Sorter100|8862_ , \new_Sorter100|8863_ , \new_Sorter100|8864_ ,
    \new_Sorter100|8865_ , \new_Sorter100|8866_ , \new_Sorter100|8867_ ,
    \new_Sorter100|8868_ , \new_Sorter100|8869_ , \new_Sorter100|8870_ ,
    \new_Sorter100|8871_ , \new_Sorter100|8872_ , \new_Sorter100|8873_ ,
    \new_Sorter100|8874_ , \new_Sorter100|8875_ , \new_Sorter100|8876_ ,
    \new_Sorter100|8877_ , \new_Sorter100|8878_ , \new_Sorter100|8879_ ,
    \new_Sorter100|8880_ , \new_Sorter100|8881_ , \new_Sorter100|8882_ ,
    \new_Sorter100|8883_ , \new_Sorter100|8884_ , \new_Sorter100|8885_ ,
    \new_Sorter100|8886_ , \new_Sorter100|8887_ , \new_Sorter100|8888_ ,
    \new_Sorter100|8889_ , \new_Sorter100|8890_ , \new_Sorter100|8891_ ,
    \new_Sorter100|8892_ , \new_Sorter100|8893_ , \new_Sorter100|8894_ ,
    \new_Sorter100|8895_ , \new_Sorter100|8896_ , \new_Sorter100|8897_ ,
    \new_Sorter100|8898_ , \new_Sorter100|8899_ , \new_Sorter100|8900_ ,
    \new_Sorter100|8999_ , \new_Sorter100|8901_ , \new_Sorter100|8902_ ,
    \new_Sorter100|8903_ , \new_Sorter100|8904_ , \new_Sorter100|8905_ ,
    \new_Sorter100|8906_ , \new_Sorter100|8907_ , \new_Sorter100|8908_ ,
    \new_Sorter100|8909_ , \new_Sorter100|8910_ , \new_Sorter100|8911_ ,
    \new_Sorter100|8912_ , \new_Sorter100|8913_ , \new_Sorter100|8914_ ,
    \new_Sorter100|8915_ , \new_Sorter100|8916_ , \new_Sorter100|8917_ ,
    \new_Sorter100|8918_ , \new_Sorter100|8919_ , \new_Sorter100|8920_ ,
    \new_Sorter100|8921_ , \new_Sorter100|8922_ , \new_Sorter100|8923_ ,
    \new_Sorter100|8924_ , \new_Sorter100|8925_ , \new_Sorter100|8926_ ,
    \new_Sorter100|8927_ , \new_Sorter100|8928_ , \new_Sorter100|8929_ ,
    \new_Sorter100|8930_ , \new_Sorter100|8931_ , \new_Sorter100|8932_ ,
    \new_Sorter100|8933_ , \new_Sorter100|8934_ , \new_Sorter100|8935_ ,
    \new_Sorter100|8936_ , \new_Sorter100|8937_ , \new_Sorter100|8938_ ,
    \new_Sorter100|8939_ , \new_Sorter100|8940_ , \new_Sorter100|8941_ ,
    \new_Sorter100|8942_ , \new_Sorter100|8943_ , \new_Sorter100|8944_ ,
    \new_Sorter100|8945_ , \new_Sorter100|8946_ , \new_Sorter100|8947_ ,
    \new_Sorter100|8948_ , \new_Sorter100|8949_ , \new_Sorter100|8950_ ,
    \new_Sorter100|8951_ , \new_Sorter100|8952_ , \new_Sorter100|8953_ ,
    \new_Sorter100|8954_ , \new_Sorter100|8955_ , \new_Sorter100|8956_ ,
    \new_Sorter100|8957_ , \new_Sorter100|8958_ , \new_Sorter100|8959_ ,
    \new_Sorter100|8960_ , \new_Sorter100|8961_ , \new_Sorter100|8962_ ,
    \new_Sorter100|8963_ , \new_Sorter100|8964_ , \new_Sorter100|8965_ ,
    \new_Sorter100|8966_ , \new_Sorter100|8967_ , \new_Sorter100|8968_ ,
    \new_Sorter100|8969_ , \new_Sorter100|8970_ , \new_Sorter100|8971_ ,
    \new_Sorter100|8972_ , \new_Sorter100|8973_ , \new_Sorter100|8974_ ,
    \new_Sorter100|8975_ , \new_Sorter100|8976_ , \new_Sorter100|8977_ ,
    \new_Sorter100|8978_ , \new_Sorter100|8979_ , \new_Sorter100|8980_ ,
    \new_Sorter100|8981_ , \new_Sorter100|8982_ , \new_Sorter100|8983_ ,
    \new_Sorter100|8984_ , \new_Sorter100|8985_ , \new_Sorter100|8986_ ,
    \new_Sorter100|8987_ , \new_Sorter100|8988_ , \new_Sorter100|8989_ ,
    \new_Sorter100|8990_ , \new_Sorter100|8991_ , \new_Sorter100|8992_ ,
    \new_Sorter100|8993_ , \new_Sorter100|8994_ , \new_Sorter100|8995_ ,
    \new_Sorter100|8996_ , \new_Sorter100|8997_ , \new_Sorter100|8998_ ,
    \new_Sorter100|9000_ , \new_Sorter100|9001_ , \new_Sorter100|9002_ ,
    \new_Sorter100|9003_ , \new_Sorter100|9004_ , \new_Sorter100|9005_ ,
    \new_Sorter100|9006_ , \new_Sorter100|9007_ , \new_Sorter100|9008_ ,
    \new_Sorter100|9009_ , \new_Sorter100|9010_ , \new_Sorter100|9011_ ,
    \new_Sorter100|9012_ , \new_Sorter100|9013_ , \new_Sorter100|9014_ ,
    \new_Sorter100|9015_ , \new_Sorter100|9016_ , \new_Sorter100|9017_ ,
    \new_Sorter100|9018_ , \new_Sorter100|9019_ , \new_Sorter100|9020_ ,
    \new_Sorter100|9021_ , \new_Sorter100|9022_ , \new_Sorter100|9023_ ,
    \new_Sorter100|9024_ , \new_Sorter100|9025_ , \new_Sorter100|9026_ ,
    \new_Sorter100|9027_ , \new_Sorter100|9028_ , \new_Sorter100|9029_ ,
    \new_Sorter100|9030_ , \new_Sorter100|9031_ , \new_Sorter100|9032_ ,
    \new_Sorter100|9033_ , \new_Sorter100|9034_ , \new_Sorter100|9035_ ,
    \new_Sorter100|9036_ , \new_Sorter100|9037_ , \new_Sorter100|9038_ ,
    \new_Sorter100|9039_ , \new_Sorter100|9040_ , \new_Sorter100|9041_ ,
    \new_Sorter100|9042_ , \new_Sorter100|9043_ , \new_Sorter100|9044_ ,
    \new_Sorter100|9045_ , \new_Sorter100|9046_ , \new_Sorter100|9047_ ,
    \new_Sorter100|9048_ , \new_Sorter100|9049_ , \new_Sorter100|9050_ ,
    \new_Sorter100|9051_ , \new_Sorter100|9052_ , \new_Sorter100|9053_ ,
    \new_Sorter100|9054_ , \new_Sorter100|9055_ , \new_Sorter100|9056_ ,
    \new_Sorter100|9057_ , \new_Sorter100|9058_ , \new_Sorter100|9059_ ,
    \new_Sorter100|9060_ , \new_Sorter100|9061_ , \new_Sorter100|9062_ ,
    \new_Sorter100|9063_ , \new_Sorter100|9064_ , \new_Sorter100|9065_ ,
    \new_Sorter100|9066_ , \new_Sorter100|9067_ , \new_Sorter100|9068_ ,
    \new_Sorter100|9069_ , \new_Sorter100|9070_ , \new_Sorter100|9071_ ,
    \new_Sorter100|9072_ , \new_Sorter100|9073_ , \new_Sorter100|9074_ ,
    \new_Sorter100|9075_ , \new_Sorter100|9076_ , \new_Sorter100|9077_ ,
    \new_Sorter100|9078_ , \new_Sorter100|9079_ , \new_Sorter100|9080_ ,
    \new_Sorter100|9081_ , \new_Sorter100|9082_ , \new_Sorter100|9083_ ,
    \new_Sorter100|9084_ , \new_Sorter100|9085_ , \new_Sorter100|9086_ ,
    \new_Sorter100|9087_ , \new_Sorter100|9088_ , \new_Sorter100|9089_ ,
    \new_Sorter100|9090_ , \new_Sorter100|9091_ , \new_Sorter100|9092_ ,
    \new_Sorter100|9093_ , \new_Sorter100|9094_ , \new_Sorter100|9095_ ,
    \new_Sorter100|9096_ , \new_Sorter100|9097_ , \new_Sorter100|9098_ ,
    \new_Sorter100|9099_ , \new_Sorter100|9100_ , \new_Sorter100|9199_ ,
    \new_Sorter100|9101_ , \new_Sorter100|9102_ , \new_Sorter100|9103_ ,
    \new_Sorter100|9104_ , \new_Sorter100|9105_ , \new_Sorter100|9106_ ,
    \new_Sorter100|9107_ , \new_Sorter100|9108_ , \new_Sorter100|9109_ ,
    \new_Sorter100|9110_ , \new_Sorter100|9111_ , \new_Sorter100|9112_ ,
    \new_Sorter100|9113_ , \new_Sorter100|9114_ , \new_Sorter100|9115_ ,
    \new_Sorter100|9116_ , \new_Sorter100|9117_ , \new_Sorter100|9118_ ,
    \new_Sorter100|9119_ , \new_Sorter100|9120_ , \new_Sorter100|9121_ ,
    \new_Sorter100|9122_ , \new_Sorter100|9123_ , \new_Sorter100|9124_ ,
    \new_Sorter100|9125_ , \new_Sorter100|9126_ , \new_Sorter100|9127_ ,
    \new_Sorter100|9128_ , \new_Sorter100|9129_ , \new_Sorter100|9130_ ,
    \new_Sorter100|9131_ , \new_Sorter100|9132_ , \new_Sorter100|9133_ ,
    \new_Sorter100|9134_ , \new_Sorter100|9135_ , \new_Sorter100|9136_ ,
    \new_Sorter100|9137_ , \new_Sorter100|9138_ , \new_Sorter100|9139_ ,
    \new_Sorter100|9140_ , \new_Sorter100|9141_ , \new_Sorter100|9142_ ,
    \new_Sorter100|9143_ , \new_Sorter100|9144_ , \new_Sorter100|9145_ ,
    \new_Sorter100|9146_ , \new_Sorter100|9147_ , \new_Sorter100|9148_ ,
    \new_Sorter100|9149_ , \new_Sorter100|9150_ , \new_Sorter100|9151_ ,
    \new_Sorter100|9152_ , \new_Sorter100|9153_ , \new_Sorter100|9154_ ,
    \new_Sorter100|9155_ , \new_Sorter100|9156_ , \new_Sorter100|9157_ ,
    \new_Sorter100|9158_ , \new_Sorter100|9159_ , \new_Sorter100|9160_ ,
    \new_Sorter100|9161_ , \new_Sorter100|9162_ , \new_Sorter100|9163_ ,
    \new_Sorter100|9164_ , \new_Sorter100|9165_ , \new_Sorter100|9166_ ,
    \new_Sorter100|9167_ , \new_Sorter100|9168_ , \new_Sorter100|9169_ ,
    \new_Sorter100|9170_ , \new_Sorter100|9171_ , \new_Sorter100|9172_ ,
    \new_Sorter100|9173_ , \new_Sorter100|9174_ , \new_Sorter100|9175_ ,
    \new_Sorter100|9176_ , \new_Sorter100|9177_ , \new_Sorter100|9178_ ,
    \new_Sorter100|9179_ , \new_Sorter100|9180_ , \new_Sorter100|9181_ ,
    \new_Sorter100|9182_ , \new_Sorter100|9183_ , \new_Sorter100|9184_ ,
    \new_Sorter100|9185_ , \new_Sorter100|9186_ , \new_Sorter100|9187_ ,
    \new_Sorter100|9188_ , \new_Sorter100|9189_ , \new_Sorter100|9190_ ,
    \new_Sorter100|9191_ , \new_Sorter100|9192_ , \new_Sorter100|9193_ ,
    \new_Sorter100|9194_ , \new_Sorter100|9195_ , \new_Sorter100|9196_ ,
    \new_Sorter100|9197_ , \new_Sorter100|9198_ , \new_Sorter100|9200_ ,
    \new_Sorter100|9201_ , \new_Sorter100|9202_ , \new_Sorter100|9203_ ,
    \new_Sorter100|9204_ , \new_Sorter100|9205_ , \new_Sorter100|9206_ ,
    \new_Sorter100|9207_ , \new_Sorter100|9208_ , \new_Sorter100|9209_ ,
    \new_Sorter100|9210_ , \new_Sorter100|9211_ , \new_Sorter100|9212_ ,
    \new_Sorter100|9213_ , \new_Sorter100|9214_ , \new_Sorter100|9215_ ,
    \new_Sorter100|9216_ , \new_Sorter100|9217_ , \new_Sorter100|9218_ ,
    \new_Sorter100|9219_ , \new_Sorter100|9220_ , \new_Sorter100|9221_ ,
    \new_Sorter100|9222_ , \new_Sorter100|9223_ , \new_Sorter100|9224_ ,
    \new_Sorter100|9225_ , \new_Sorter100|9226_ , \new_Sorter100|9227_ ,
    \new_Sorter100|9228_ , \new_Sorter100|9229_ , \new_Sorter100|9230_ ,
    \new_Sorter100|9231_ , \new_Sorter100|9232_ , \new_Sorter100|9233_ ,
    \new_Sorter100|9234_ , \new_Sorter100|9235_ , \new_Sorter100|9236_ ,
    \new_Sorter100|9237_ , \new_Sorter100|9238_ , \new_Sorter100|9239_ ,
    \new_Sorter100|9240_ , \new_Sorter100|9241_ , \new_Sorter100|9242_ ,
    \new_Sorter100|9243_ , \new_Sorter100|9244_ , \new_Sorter100|9245_ ,
    \new_Sorter100|9246_ , \new_Sorter100|9247_ , \new_Sorter100|9248_ ,
    \new_Sorter100|9249_ , \new_Sorter100|9250_ , \new_Sorter100|9251_ ,
    \new_Sorter100|9252_ , \new_Sorter100|9253_ , \new_Sorter100|9254_ ,
    \new_Sorter100|9255_ , \new_Sorter100|9256_ , \new_Sorter100|9257_ ,
    \new_Sorter100|9258_ , \new_Sorter100|9259_ , \new_Sorter100|9260_ ,
    \new_Sorter100|9261_ , \new_Sorter100|9262_ , \new_Sorter100|9263_ ,
    \new_Sorter100|9264_ , \new_Sorter100|9265_ , \new_Sorter100|9266_ ,
    \new_Sorter100|9267_ , \new_Sorter100|9268_ , \new_Sorter100|9269_ ,
    \new_Sorter100|9270_ , \new_Sorter100|9271_ , \new_Sorter100|9272_ ,
    \new_Sorter100|9273_ , \new_Sorter100|9274_ , \new_Sorter100|9275_ ,
    \new_Sorter100|9276_ , \new_Sorter100|9277_ , \new_Sorter100|9278_ ,
    \new_Sorter100|9279_ , \new_Sorter100|9280_ , \new_Sorter100|9281_ ,
    \new_Sorter100|9282_ , \new_Sorter100|9283_ , \new_Sorter100|9284_ ,
    \new_Sorter100|9285_ , \new_Sorter100|9286_ , \new_Sorter100|9287_ ,
    \new_Sorter100|9288_ , \new_Sorter100|9289_ , \new_Sorter100|9290_ ,
    \new_Sorter100|9291_ , \new_Sorter100|9292_ , \new_Sorter100|9293_ ,
    \new_Sorter100|9294_ , \new_Sorter100|9295_ , \new_Sorter100|9296_ ,
    \new_Sorter100|9297_ , \new_Sorter100|9298_ , \new_Sorter100|9299_ ,
    \new_Sorter100|9300_ , \new_Sorter100|9399_ , \new_Sorter100|9301_ ,
    \new_Sorter100|9302_ , \new_Sorter100|9303_ , \new_Sorter100|9304_ ,
    \new_Sorter100|9305_ , \new_Sorter100|9306_ , \new_Sorter100|9307_ ,
    \new_Sorter100|9308_ , \new_Sorter100|9309_ , \new_Sorter100|9310_ ,
    \new_Sorter100|9311_ , \new_Sorter100|9312_ , \new_Sorter100|9313_ ,
    \new_Sorter100|9314_ , \new_Sorter100|9315_ , \new_Sorter100|9316_ ,
    \new_Sorter100|9317_ , \new_Sorter100|9318_ , \new_Sorter100|9319_ ,
    \new_Sorter100|9320_ , \new_Sorter100|9321_ , \new_Sorter100|9322_ ,
    \new_Sorter100|9323_ , \new_Sorter100|9324_ , \new_Sorter100|9325_ ,
    \new_Sorter100|9326_ , \new_Sorter100|9327_ , \new_Sorter100|9328_ ,
    \new_Sorter100|9329_ , \new_Sorter100|9330_ , \new_Sorter100|9331_ ,
    \new_Sorter100|9332_ , \new_Sorter100|9333_ , \new_Sorter100|9334_ ,
    \new_Sorter100|9335_ , \new_Sorter100|9336_ , \new_Sorter100|9337_ ,
    \new_Sorter100|9338_ , \new_Sorter100|9339_ , \new_Sorter100|9340_ ,
    \new_Sorter100|9341_ , \new_Sorter100|9342_ , \new_Sorter100|9343_ ,
    \new_Sorter100|9344_ , \new_Sorter100|9345_ , \new_Sorter100|9346_ ,
    \new_Sorter100|9347_ , \new_Sorter100|9348_ , \new_Sorter100|9349_ ,
    \new_Sorter100|9350_ , \new_Sorter100|9351_ , \new_Sorter100|9352_ ,
    \new_Sorter100|9353_ , \new_Sorter100|9354_ , \new_Sorter100|9355_ ,
    \new_Sorter100|9356_ , \new_Sorter100|9357_ , \new_Sorter100|9358_ ,
    \new_Sorter100|9359_ , \new_Sorter100|9360_ , \new_Sorter100|9361_ ,
    \new_Sorter100|9362_ , \new_Sorter100|9363_ , \new_Sorter100|9364_ ,
    \new_Sorter100|9365_ , \new_Sorter100|9366_ , \new_Sorter100|9367_ ,
    \new_Sorter100|9368_ , \new_Sorter100|9369_ , \new_Sorter100|9370_ ,
    \new_Sorter100|9371_ , \new_Sorter100|9372_ , \new_Sorter100|9373_ ,
    \new_Sorter100|9374_ , \new_Sorter100|9375_ , \new_Sorter100|9376_ ,
    \new_Sorter100|9377_ , \new_Sorter100|9378_ , \new_Sorter100|9379_ ,
    \new_Sorter100|9380_ , \new_Sorter100|9381_ , \new_Sorter100|9382_ ,
    \new_Sorter100|9383_ , \new_Sorter100|9384_ , \new_Sorter100|9385_ ,
    \new_Sorter100|9386_ , \new_Sorter100|9387_ , \new_Sorter100|9388_ ,
    \new_Sorter100|9389_ , \new_Sorter100|9390_ , \new_Sorter100|9391_ ,
    \new_Sorter100|9392_ , \new_Sorter100|9393_ , \new_Sorter100|9394_ ,
    \new_Sorter100|9395_ , \new_Sorter100|9396_ , \new_Sorter100|9397_ ,
    \new_Sorter100|9398_ , \new_Sorter100|9400_ , \new_Sorter100|9401_ ,
    \new_Sorter100|9402_ , \new_Sorter100|9403_ , \new_Sorter100|9404_ ,
    \new_Sorter100|9405_ , \new_Sorter100|9406_ , \new_Sorter100|9407_ ,
    \new_Sorter100|9408_ , \new_Sorter100|9409_ , \new_Sorter100|9410_ ,
    \new_Sorter100|9411_ , \new_Sorter100|9412_ , \new_Sorter100|9413_ ,
    \new_Sorter100|9414_ , \new_Sorter100|9415_ , \new_Sorter100|9416_ ,
    \new_Sorter100|9417_ , \new_Sorter100|9418_ , \new_Sorter100|9419_ ,
    \new_Sorter100|9420_ , \new_Sorter100|9421_ , \new_Sorter100|9422_ ,
    \new_Sorter100|9423_ , \new_Sorter100|9424_ , \new_Sorter100|9425_ ,
    \new_Sorter100|9426_ , \new_Sorter100|9427_ , \new_Sorter100|9428_ ,
    \new_Sorter100|9429_ , \new_Sorter100|9430_ , \new_Sorter100|9431_ ,
    \new_Sorter100|9432_ , \new_Sorter100|9433_ , \new_Sorter100|9434_ ,
    \new_Sorter100|9435_ , \new_Sorter100|9436_ , \new_Sorter100|9437_ ,
    \new_Sorter100|9438_ , \new_Sorter100|9439_ , \new_Sorter100|9440_ ,
    \new_Sorter100|9441_ , \new_Sorter100|9442_ , \new_Sorter100|9443_ ,
    \new_Sorter100|9444_ , \new_Sorter100|9445_ , \new_Sorter100|9446_ ,
    \new_Sorter100|9447_ , \new_Sorter100|9448_ , \new_Sorter100|9449_ ,
    \new_Sorter100|9450_ , \new_Sorter100|9451_ , \new_Sorter100|9452_ ,
    \new_Sorter100|9453_ , \new_Sorter100|9454_ , \new_Sorter100|9455_ ,
    \new_Sorter100|9456_ , \new_Sorter100|9457_ , \new_Sorter100|9458_ ,
    \new_Sorter100|9459_ , \new_Sorter100|9460_ , \new_Sorter100|9461_ ,
    \new_Sorter100|9462_ , \new_Sorter100|9463_ , \new_Sorter100|9464_ ,
    \new_Sorter100|9465_ , \new_Sorter100|9466_ , \new_Sorter100|9467_ ,
    \new_Sorter100|9468_ , \new_Sorter100|9469_ , \new_Sorter100|9470_ ,
    \new_Sorter100|9471_ , \new_Sorter100|9472_ , \new_Sorter100|9473_ ,
    \new_Sorter100|9474_ , \new_Sorter100|9475_ , \new_Sorter100|9476_ ,
    \new_Sorter100|9477_ , \new_Sorter100|9478_ , \new_Sorter100|9479_ ,
    \new_Sorter100|9480_ , \new_Sorter100|9481_ , \new_Sorter100|9482_ ,
    \new_Sorter100|9483_ , \new_Sorter100|9484_ , \new_Sorter100|9485_ ,
    \new_Sorter100|9486_ , \new_Sorter100|9487_ , \new_Sorter100|9488_ ,
    \new_Sorter100|9489_ , \new_Sorter100|9490_ , \new_Sorter100|9491_ ,
    \new_Sorter100|9492_ , \new_Sorter100|9493_ , \new_Sorter100|9494_ ,
    \new_Sorter100|9495_ , \new_Sorter100|9496_ , \new_Sorter100|9497_ ,
    \new_Sorter100|9498_ , \new_Sorter100|9499_ , \new_Sorter100|9500_ ,
    \new_Sorter100|9599_ , \new_Sorter100|9501_ , \new_Sorter100|9502_ ,
    \new_Sorter100|9503_ , \new_Sorter100|9504_ , \new_Sorter100|9505_ ,
    \new_Sorter100|9506_ , \new_Sorter100|9507_ , \new_Sorter100|9508_ ,
    \new_Sorter100|9509_ , \new_Sorter100|9510_ , \new_Sorter100|9511_ ,
    \new_Sorter100|9512_ , \new_Sorter100|9513_ , \new_Sorter100|9514_ ,
    \new_Sorter100|9515_ , \new_Sorter100|9516_ , \new_Sorter100|9517_ ,
    \new_Sorter100|9518_ , \new_Sorter100|9519_ , \new_Sorter100|9520_ ,
    \new_Sorter100|9521_ , \new_Sorter100|9522_ , \new_Sorter100|9523_ ,
    \new_Sorter100|9524_ , \new_Sorter100|9525_ , \new_Sorter100|9526_ ,
    \new_Sorter100|9527_ , \new_Sorter100|9528_ , \new_Sorter100|9529_ ,
    \new_Sorter100|9530_ , \new_Sorter100|9531_ , \new_Sorter100|9532_ ,
    \new_Sorter100|9533_ , \new_Sorter100|9534_ , \new_Sorter100|9535_ ,
    \new_Sorter100|9536_ , \new_Sorter100|9537_ , \new_Sorter100|9538_ ,
    \new_Sorter100|9539_ , \new_Sorter100|9540_ , \new_Sorter100|9541_ ,
    \new_Sorter100|9542_ , \new_Sorter100|9543_ , \new_Sorter100|9544_ ,
    \new_Sorter100|9545_ , \new_Sorter100|9546_ , \new_Sorter100|9547_ ,
    \new_Sorter100|9548_ , \new_Sorter100|9549_ , \new_Sorter100|9550_ ,
    \new_Sorter100|9551_ , \new_Sorter100|9552_ , \new_Sorter100|9553_ ,
    \new_Sorter100|9554_ , \new_Sorter100|9555_ , \new_Sorter100|9556_ ,
    \new_Sorter100|9557_ , \new_Sorter100|9558_ , \new_Sorter100|9559_ ,
    \new_Sorter100|9560_ , \new_Sorter100|9561_ , \new_Sorter100|9562_ ,
    \new_Sorter100|9563_ , \new_Sorter100|9564_ , \new_Sorter100|9565_ ,
    \new_Sorter100|9566_ , \new_Sorter100|9567_ , \new_Sorter100|9568_ ,
    \new_Sorter100|9569_ , \new_Sorter100|9570_ , \new_Sorter100|9571_ ,
    \new_Sorter100|9572_ , \new_Sorter100|9573_ , \new_Sorter100|9574_ ,
    \new_Sorter100|9575_ , \new_Sorter100|9576_ , \new_Sorter100|9577_ ,
    \new_Sorter100|9578_ , \new_Sorter100|9579_ , \new_Sorter100|9580_ ,
    \new_Sorter100|9581_ , \new_Sorter100|9582_ , \new_Sorter100|9583_ ,
    \new_Sorter100|9584_ , \new_Sorter100|9585_ , \new_Sorter100|9586_ ,
    \new_Sorter100|9587_ , \new_Sorter100|9588_ , \new_Sorter100|9589_ ,
    \new_Sorter100|9590_ , \new_Sorter100|9591_ , \new_Sorter100|9592_ ,
    \new_Sorter100|9593_ , \new_Sorter100|9594_ , \new_Sorter100|9595_ ,
    \new_Sorter100|9596_ , \new_Sorter100|9597_ , \new_Sorter100|9598_ ,
    \new_Sorter100|9600_ , \new_Sorter100|9601_ , \new_Sorter100|9602_ ,
    \new_Sorter100|9603_ , \new_Sorter100|9604_ , \new_Sorter100|9605_ ,
    \new_Sorter100|9606_ , \new_Sorter100|9607_ , \new_Sorter100|9608_ ,
    \new_Sorter100|9609_ , \new_Sorter100|9610_ , \new_Sorter100|9611_ ,
    \new_Sorter100|9612_ , \new_Sorter100|9613_ , \new_Sorter100|9614_ ,
    \new_Sorter100|9615_ , \new_Sorter100|9616_ , \new_Sorter100|9617_ ,
    \new_Sorter100|9618_ , \new_Sorter100|9619_ , \new_Sorter100|9620_ ,
    \new_Sorter100|9621_ , \new_Sorter100|9622_ , \new_Sorter100|9623_ ,
    \new_Sorter100|9624_ , \new_Sorter100|9625_ , \new_Sorter100|9626_ ,
    \new_Sorter100|9627_ , \new_Sorter100|9628_ , \new_Sorter100|9629_ ,
    \new_Sorter100|9630_ , \new_Sorter100|9631_ , \new_Sorter100|9632_ ,
    \new_Sorter100|9633_ , \new_Sorter100|9634_ , \new_Sorter100|9635_ ,
    \new_Sorter100|9636_ , \new_Sorter100|9637_ , \new_Sorter100|9638_ ,
    \new_Sorter100|9639_ , \new_Sorter100|9640_ , \new_Sorter100|9641_ ,
    \new_Sorter100|9642_ , \new_Sorter100|9643_ , \new_Sorter100|9644_ ,
    \new_Sorter100|9645_ , \new_Sorter100|9646_ , \new_Sorter100|9647_ ,
    \new_Sorter100|9648_ , \new_Sorter100|9649_ , \new_Sorter100|9650_ ,
    \new_Sorter100|9651_ , \new_Sorter100|9652_ , \new_Sorter100|9653_ ,
    \new_Sorter100|9654_ , \new_Sorter100|9655_ , \new_Sorter100|9656_ ,
    \new_Sorter100|9657_ , \new_Sorter100|9658_ , \new_Sorter100|9659_ ,
    \new_Sorter100|9660_ , \new_Sorter100|9661_ , \new_Sorter100|9662_ ,
    \new_Sorter100|9663_ , \new_Sorter100|9664_ , \new_Sorter100|9665_ ,
    \new_Sorter100|9666_ , \new_Sorter100|9667_ , \new_Sorter100|9668_ ,
    \new_Sorter100|9669_ , \new_Sorter100|9670_ , \new_Sorter100|9671_ ,
    \new_Sorter100|9672_ , \new_Sorter100|9673_ , \new_Sorter100|9674_ ,
    \new_Sorter100|9675_ , \new_Sorter100|9676_ , \new_Sorter100|9677_ ,
    \new_Sorter100|9678_ , \new_Sorter100|9679_ , \new_Sorter100|9680_ ,
    \new_Sorter100|9681_ , \new_Sorter100|9682_ , \new_Sorter100|9683_ ,
    \new_Sorter100|9684_ , \new_Sorter100|9685_ , \new_Sorter100|9686_ ,
    \new_Sorter100|9687_ , \new_Sorter100|9688_ , \new_Sorter100|9689_ ,
    \new_Sorter100|9690_ , \new_Sorter100|9691_ , \new_Sorter100|9692_ ,
    \new_Sorter100|9693_ , \new_Sorter100|9694_ , \new_Sorter100|9695_ ,
    \new_Sorter100|9696_ , \new_Sorter100|9697_ , \new_Sorter100|9698_ ,
    \new_Sorter100|9699_ , \new_Sorter100|9700_ , \new_Sorter100|9799_ ,
    \new_Sorter100|9701_ , \new_Sorter100|9702_ , \new_Sorter100|9703_ ,
    \new_Sorter100|9704_ , \new_Sorter100|9705_ , \new_Sorter100|9706_ ,
    \new_Sorter100|9707_ , \new_Sorter100|9708_ , \new_Sorter100|9709_ ,
    \new_Sorter100|9710_ , \new_Sorter100|9711_ , \new_Sorter100|9712_ ,
    \new_Sorter100|9713_ , \new_Sorter100|9714_ , \new_Sorter100|9715_ ,
    \new_Sorter100|9716_ , \new_Sorter100|9717_ , \new_Sorter100|9718_ ,
    \new_Sorter100|9719_ , \new_Sorter100|9720_ , \new_Sorter100|9721_ ,
    \new_Sorter100|9722_ , \new_Sorter100|9723_ , \new_Sorter100|9724_ ,
    \new_Sorter100|9725_ , \new_Sorter100|9726_ , \new_Sorter100|9727_ ,
    \new_Sorter100|9728_ , \new_Sorter100|9729_ , \new_Sorter100|9730_ ,
    \new_Sorter100|9731_ , \new_Sorter100|9732_ , \new_Sorter100|9733_ ,
    \new_Sorter100|9734_ , \new_Sorter100|9735_ , \new_Sorter100|9736_ ,
    \new_Sorter100|9737_ , \new_Sorter100|9738_ , \new_Sorter100|9739_ ,
    \new_Sorter100|9740_ , \new_Sorter100|9741_ , \new_Sorter100|9742_ ,
    \new_Sorter100|9743_ , \new_Sorter100|9744_ , \new_Sorter100|9745_ ,
    \new_Sorter100|9746_ , \new_Sorter100|9747_ , \new_Sorter100|9748_ ,
    \new_Sorter100|9749_ , \new_Sorter100|9750_ , \new_Sorter100|9751_ ,
    \new_Sorter100|9752_ , \new_Sorter100|9753_ , \new_Sorter100|9754_ ,
    \new_Sorter100|9755_ , \new_Sorter100|9756_ , \new_Sorter100|9757_ ,
    \new_Sorter100|9758_ , \new_Sorter100|9759_ , \new_Sorter100|9760_ ,
    \new_Sorter100|9761_ , \new_Sorter100|9762_ , \new_Sorter100|9763_ ,
    \new_Sorter100|9764_ , \new_Sorter100|9765_ , \new_Sorter100|9766_ ,
    \new_Sorter100|9767_ , \new_Sorter100|9768_ , \new_Sorter100|9769_ ,
    \new_Sorter100|9770_ , \new_Sorter100|9771_ , \new_Sorter100|9772_ ,
    \new_Sorter100|9773_ , \new_Sorter100|9774_ , \new_Sorter100|9775_ ,
    \new_Sorter100|9776_ , \new_Sorter100|9777_ , \new_Sorter100|9778_ ,
    \new_Sorter100|9779_ , \new_Sorter100|9780_ , \new_Sorter100|9781_ ,
    \new_Sorter100|9782_ , \new_Sorter100|9783_ , \new_Sorter100|9784_ ,
    \new_Sorter100|9785_ , \new_Sorter100|9786_ , \new_Sorter100|9787_ ,
    \new_Sorter100|9788_ , \new_Sorter100|9789_ , \new_Sorter100|9790_ ,
    \new_Sorter100|9791_ , \new_Sorter100|9792_ , \new_Sorter100|9793_ ,
    \new_Sorter100|9794_ , \new_Sorter100|9795_ , \new_Sorter100|9796_ ,
    \new_Sorter100|9797_ , \new_Sorter100|9798_ , \new_Sorter100|9800_ ,
    \new_Sorter100|9801_ , \new_Sorter100|9802_ , \new_Sorter100|9803_ ,
    \new_Sorter100|9804_ , \new_Sorter100|9805_ , \new_Sorter100|9806_ ,
    \new_Sorter100|9807_ , \new_Sorter100|9808_ , \new_Sorter100|9809_ ,
    \new_Sorter100|9810_ , \new_Sorter100|9811_ , \new_Sorter100|9812_ ,
    \new_Sorter100|9813_ , \new_Sorter100|9814_ , \new_Sorter100|9815_ ,
    \new_Sorter100|9816_ , \new_Sorter100|9817_ , \new_Sorter100|9818_ ,
    \new_Sorter100|9819_ , \new_Sorter100|9820_ , \new_Sorter100|9821_ ,
    \new_Sorter100|9822_ , \new_Sorter100|9823_ , \new_Sorter100|9824_ ,
    \new_Sorter100|9825_ , \new_Sorter100|9826_ , \new_Sorter100|9827_ ,
    \new_Sorter100|9828_ , \new_Sorter100|9829_ , \new_Sorter100|9830_ ,
    \new_Sorter100|9831_ , \new_Sorter100|9832_ , \new_Sorter100|9833_ ,
    \new_Sorter100|9834_ , \new_Sorter100|9835_ , \new_Sorter100|9836_ ,
    \new_Sorter100|9837_ , \new_Sorter100|9838_ , \new_Sorter100|9839_ ,
    \new_Sorter100|9840_ , \new_Sorter100|9841_ , \new_Sorter100|9842_ ,
    \new_Sorter100|9843_ , \new_Sorter100|9844_ , \new_Sorter100|9845_ ,
    \new_Sorter100|9846_ , \new_Sorter100|9847_ , \new_Sorter100|9848_ ,
    \new_Sorter100|9849_ , \new_Sorter100|9850_ , \new_Sorter100|9851_ ,
    \new_Sorter100|9852_ , \new_Sorter100|9853_ , \new_Sorter100|9854_ ,
    \new_Sorter100|9855_ , \new_Sorter100|9856_ , \new_Sorter100|9857_ ,
    \new_Sorter100|9858_ , \new_Sorter100|9859_ , \new_Sorter100|9860_ ,
    \new_Sorter100|9861_ , \new_Sorter100|9862_ , \new_Sorter100|9863_ ,
    \new_Sorter100|9864_ , \new_Sorter100|9865_ , \new_Sorter100|9866_ ,
    \new_Sorter100|9867_ , \new_Sorter100|9868_ , \new_Sorter100|9869_ ,
    \new_Sorter100|9870_ , \new_Sorter100|9871_ , \new_Sorter100|9872_ ,
    \new_Sorter100|9873_ , \new_Sorter100|9874_ , \new_Sorter100|9875_ ,
    \new_Sorter100|9876_ , \new_Sorter100|9877_ , \new_Sorter100|9878_ ,
    \new_Sorter100|9879_ , \new_Sorter100|9880_ , \new_Sorter100|9881_ ,
    \new_Sorter100|9882_ , \new_Sorter100|9883_ , \new_Sorter100|9884_ ,
    \new_Sorter100|9885_ , \new_Sorter100|9886_ , \new_Sorter100|9887_ ,
    \new_Sorter100|9888_ , \new_Sorter100|9889_ , \new_Sorter100|9890_ ,
    \new_Sorter100|9891_ , \new_Sorter100|9892_ , \new_Sorter100|9893_ ,
    \new_Sorter100|9894_ , \new_Sorter100|9895_ , \new_Sorter100|9896_ ,
    \new_Sorter100|9897_ , \new_Sorter100|9898_ , \new_Sorter100|9899_ ,
    \new_Sorter100|9900_ , \new_Sorter100|9999_ , \new_Sorter100|9901_ ,
    \new_Sorter100|9902_ , \new_Sorter100|9903_ , \new_Sorter100|9904_ ,
    \new_Sorter100|9905_ , \new_Sorter100|9906_ , \new_Sorter100|9907_ ,
    \new_Sorter100|9908_ , \new_Sorter100|9909_ , \new_Sorter100|9910_ ,
    \new_Sorter100|9911_ , \new_Sorter100|9912_ , \new_Sorter100|9913_ ,
    \new_Sorter100|9914_ , \new_Sorter100|9915_ , \new_Sorter100|9916_ ,
    \new_Sorter100|9917_ , \new_Sorter100|9918_ , \new_Sorter100|9919_ ,
    \new_Sorter100|9920_ , \new_Sorter100|9921_ , \new_Sorter100|9922_ ,
    \new_Sorter100|9923_ , \new_Sorter100|9924_ , \new_Sorter100|9925_ ,
    \new_Sorter100|9926_ , \new_Sorter100|9927_ , \new_Sorter100|9928_ ,
    \new_Sorter100|9929_ , \new_Sorter100|9930_ , \new_Sorter100|9931_ ,
    \new_Sorter100|9932_ , \new_Sorter100|9933_ , \new_Sorter100|9934_ ,
    \new_Sorter100|9935_ , \new_Sorter100|9936_ , \new_Sorter100|9937_ ,
    \new_Sorter100|9938_ , \new_Sorter100|9939_ , \new_Sorter100|9940_ ,
    \new_Sorter100|9941_ , \new_Sorter100|9942_ , \new_Sorter100|9943_ ,
    \new_Sorter100|9944_ , \new_Sorter100|9945_ , \new_Sorter100|9946_ ,
    \new_Sorter100|9947_ , \new_Sorter100|9948_ , \new_Sorter100|9949_ ,
    \new_Sorter100|9950_ , \new_Sorter100|9951_ , \new_Sorter100|9952_ ,
    \new_Sorter100|9953_ , \new_Sorter100|9954_ , \new_Sorter100|9955_ ,
    \new_Sorter100|9956_ , \new_Sorter100|9957_ , \new_Sorter100|9958_ ,
    \new_Sorter100|9959_ , \new_Sorter100|9960_ , \new_Sorter100|9961_ ,
    \new_Sorter100|9962_ , \new_Sorter100|9963_ , \new_Sorter100|9964_ ,
    \new_Sorter100|9965_ , \new_Sorter100|9966_ , \new_Sorter100|9967_ ,
    \new_Sorter100|9968_ , \new_Sorter100|9969_ , \new_Sorter100|9970_ ,
    \new_Sorter100|9971_ , \new_Sorter100|9972_ , \new_Sorter100|9973_ ,
    \new_Sorter100|9974_ , \new_Sorter100|9975_ , \new_Sorter100|9976_ ,
    \new_Sorter100|9977_ , \new_Sorter100|9978_ , \new_Sorter100|9979_ ,
    \new_Sorter100|9980_ , \new_Sorter100|9981_ , \new_Sorter100|9982_ ,
    \new_Sorter100|9983_ , \new_Sorter100|9984_ , \new_Sorter100|9985_ ,
    \new_Sorter100|9986_ , \new_Sorter100|9987_ , \new_Sorter100|9988_ ,
    \new_Sorter100|9989_ , \new_Sorter100|9990_ , \new_Sorter100|9991_ ,
    \new_Sorter100|9992_ , \new_Sorter100|9993_ , \new_Sorter100|9994_ ,
    \new_Sorter100|9995_ , \new_Sorter100|9996_ , \new_Sorter100|9997_ ,
    \new_Sorter100|9998_ , \new_Sorter100|10000_ , \new_Sorter100|10001_ ,
    \new_Sorter100|10002_ , \new_Sorter100|10003_ , \new_Sorter100|10004_ ,
    \new_Sorter100|10005_ , \new_Sorter100|10006_ , \new_Sorter100|10007_ ,
    \new_Sorter100|10008_ , \new_Sorter100|10009_ , \new_Sorter100|10010_ ,
    \new_Sorter100|10011_ , \new_Sorter100|10012_ , \new_Sorter100|10013_ ,
    \new_Sorter100|10014_ , \new_Sorter100|10015_ , \new_Sorter100|10016_ ,
    \new_Sorter100|10017_ , \new_Sorter100|10018_ , \new_Sorter100|10019_ ,
    \new_Sorter100|10020_ , \new_Sorter100|10021_ , \new_Sorter100|10022_ ,
    \new_Sorter100|10023_ , \new_Sorter100|10024_ , \new_Sorter100|10025_ ,
    \new_Sorter100|10026_ , \new_Sorter100|10027_ , \new_Sorter100|10028_ ,
    \new_Sorter100|10029_ , \new_Sorter100|10030_ , \new_Sorter100|10031_ ,
    \new_Sorter100|10032_ , \new_Sorter100|10033_ , \new_Sorter100|10034_ ,
    \new_Sorter100|10035_ , \new_Sorter100|10036_ , \new_Sorter100|10037_ ,
    \new_Sorter100|10038_ , \new_Sorter100|10039_ , \new_Sorter100|10040_ ,
    \new_Sorter100|10041_ , \new_Sorter100|10042_ , \new_Sorter100|10043_ ,
    \new_Sorter100|10044_ , \new_Sorter100|10045_ , \new_Sorter100|10046_ ,
    \new_Sorter100|10047_ , \new_Sorter100|10048_ , \new_Sorter100|10049_ ,
    \new_Sorter100|10050_ , \new_Sorter100|10051_ , \new_Sorter100|10052_ ,
    \new_Sorter100|10053_ , \new_Sorter100|10054_ , \new_Sorter100|10055_ ,
    \new_Sorter100|10056_ , \new_Sorter100|10057_ , \new_Sorter100|10058_ ,
    \new_Sorter100|10059_ , \new_Sorter100|10060_ , \new_Sorter100|10061_ ,
    \new_Sorter100|10062_ , \new_Sorter100|10063_ , \new_Sorter100|10064_ ,
    \new_Sorter100|10065_ , \new_Sorter100|10066_ , \new_Sorter100|10067_ ,
    \new_Sorter100|10068_ , \new_Sorter100|10069_ , \new_Sorter100|10070_ ,
    \new_Sorter100|10071_ , \new_Sorter100|10072_ , \new_Sorter100|10073_ ,
    \new_Sorter100|10074_ , \new_Sorter100|10075_ , \new_Sorter100|10076_ ,
    \new_Sorter100|10077_ , \new_Sorter100|10078_ , \new_Sorter100|10079_ ,
    \new_Sorter100|10080_ , \new_Sorter100|10081_ , \new_Sorter100|10082_ ,
    \new_Sorter100|10083_ , \new_Sorter100|10084_ , \new_Sorter100|10085_ ,
    \new_Sorter100|10086_ , \new_Sorter100|10087_ , \new_Sorter100|10088_ ,
    \new_Sorter100|10089_ , \new_Sorter100|10090_ , \new_Sorter100|10091_ ,
    \new_Sorter100|10092_ , \new_Sorter100|10093_ , \new_Sorter100|10094_ ,
    \new_Sorter100|10095_ , \new_Sorter100|10096_ , \new_Sorter100|10097_ ,
    \new_Sorter100|10098_ , \new_Sorter100|10099_ , \new_Sorter100|10100_ ,
    \new_Sorter100|10199_ , \new_Sorter100|10101_ , \new_Sorter100|10102_ ,
    \new_Sorter100|10103_ , \new_Sorter100|10104_ , \new_Sorter100|10105_ ,
    \new_Sorter100|10106_ , \new_Sorter100|10107_ , \new_Sorter100|10108_ ,
    \new_Sorter100|10109_ , \new_Sorter100|10110_ , \new_Sorter100|10111_ ,
    \new_Sorter100|10112_ , \new_Sorter100|10113_ , \new_Sorter100|10114_ ,
    \new_Sorter100|10115_ , \new_Sorter100|10116_ , \new_Sorter100|10117_ ,
    \new_Sorter100|10118_ , \new_Sorter100|10119_ , \new_Sorter100|10120_ ,
    \new_Sorter100|10121_ , \new_Sorter100|10122_ , \new_Sorter100|10123_ ,
    \new_Sorter100|10124_ , \new_Sorter100|10125_ , \new_Sorter100|10126_ ,
    \new_Sorter100|10127_ , \new_Sorter100|10128_ , \new_Sorter100|10129_ ,
    \new_Sorter100|10130_ , \new_Sorter100|10131_ , \new_Sorter100|10132_ ,
    \new_Sorter100|10133_ , \new_Sorter100|10134_ , \new_Sorter100|10135_ ,
    \new_Sorter100|10136_ , \new_Sorter100|10137_ , \new_Sorter100|10138_ ,
    \new_Sorter100|10139_ , \new_Sorter100|10140_ , \new_Sorter100|10141_ ,
    \new_Sorter100|10142_ , \new_Sorter100|10143_ , \new_Sorter100|10144_ ,
    \new_Sorter100|10145_ , \new_Sorter100|10146_ , \new_Sorter100|10147_ ,
    \new_Sorter100|10148_ , \new_Sorter100|10149_ , \new_Sorter100|10150_ ,
    \new_Sorter100|10151_ , \new_Sorter100|10152_ , \new_Sorter100|10153_ ,
    \new_Sorter100|10154_ , \new_Sorter100|10155_ , \new_Sorter100|10156_ ,
    \new_Sorter100|10157_ , \new_Sorter100|10158_ , \new_Sorter100|10159_ ,
    \new_Sorter100|10160_ , \new_Sorter100|10161_ , \new_Sorter100|10162_ ,
    \new_Sorter100|10163_ , \new_Sorter100|10164_ , \new_Sorter100|10165_ ,
    \new_Sorter100|10166_ , \new_Sorter100|10167_ , \new_Sorter100|10168_ ,
    \new_Sorter100|10169_ , \new_Sorter100|10170_ , \new_Sorter100|10171_ ,
    \new_Sorter100|10172_ , \new_Sorter100|10173_ , \new_Sorter100|10174_ ,
    \new_Sorter100|10175_ , \new_Sorter100|10176_ , \new_Sorter100|10177_ ,
    \new_Sorter100|10178_ , \new_Sorter100|10179_ , \new_Sorter100|10180_ ,
    \new_Sorter100|10181_ , \new_Sorter100|10182_ , \new_Sorter100|10183_ ,
    \new_Sorter100|10184_ , \new_Sorter100|10185_ , \new_Sorter100|10186_ ,
    \new_Sorter100|10187_ , \new_Sorter100|10188_ , \new_Sorter100|10189_ ,
    \new_Sorter100|10190_ , \new_Sorter100|10191_ , \new_Sorter100|10192_ ,
    \new_Sorter100|10193_ , \new_Sorter100|10194_ , \new_Sorter100|10195_ ,
    \new_Sorter100|10196_ , \new_Sorter100|10197_ , \new_Sorter100|10198_ ,
    \new_Sorter100|10200_ , \new_Sorter100|10201_ , \new_Sorter100|10202_ ,
    \new_Sorter100|10203_ , \new_Sorter100|10204_ , \new_Sorter100|10205_ ,
    \new_Sorter100|10206_ , \new_Sorter100|10207_ , \new_Sorter100|10208_ ,
    \new_Sorter100|10209_ , \new_Sorter100|10210_ , \new_Sorter100|10211_ ,
    \new_Sorter100|10212_ , \new_Sorter100|10213_ , \new_Sorter100|10214_ ,
    \new_Sorter100|10215_ , \new_Sorter100|10216_ , \new_Sorter100|10217_ ,
    \new_Sorter100|10218_ , \new_Sorter100|10219_ , \new_Sorter100|10220_ ,
    \new_Sorter100|10221_ , \new_Sorter100|10222_ , \new_Sorter100|10223_ ,
    \new_Sorter100|10224_ , \new_Sorter100|10225_ , \new_Sorter100|10226_ ,
    \new_Sorter100|10227_ , \new_Sorter100|10228_ , \new_Sorter100|10229_ ,
    \new_Sorter100|10230_ , \new_Sorter100|10231_ , \new_Sorter100|10232_ ,
    \new_Sorter100|10233_ , \new_Sorter100|10234_ , \new_Sorter100|10235_ ,
    \new_Sorter100|10236_ , \new_Sorter100|10237_ , \new_Sorter100|10238_ ,
    \new_Sorter100|10239_ , \new_Sorter100|10240_ , \new_Sorter100|10241_ ,
    \new_Sorter100|10242_ , \new_Sorter100|10243_ , \new_Sorter100|10244_ ,
    \new_Sorter100|10245_ , \new_Sorter100|10246_ , \new_Sorter100|10247_ ,
    \new_Sorter100|10248_ , \new_Sorter100|10249_ , \new_Sorter100|10250_ ,
    \new_Sorter100|10251_ , \new_Sorter100|10252_ , \new_Sorter100|10253_ ,
    \new_Sorter100|10254_ , \new_Sorter100|10255_ , \new_Sorter100|10256_ ,
    \new_Sorter100|10257_ , \new_Sorter100|10258_ , \new_Sorter100|10259_ ,
    \new_Sorter100|10260_ , \new_Sorter100|10261_ , \new_Sorter100|10262_ ,
    \new_Sorter100|10263_ , \new_Sorter100|10264_ , \new_Sorter100|10265_ ,
    \new_Sorter100|10266_ , \new_Sorter100|10267_ , \new_Sorter100|10268_ ,
    \new_Sorter100|10269_ , \new_Sorter100|10270_ , \new_Sorter100|10271_ ,
    \new_Sorter100|10272_ , \new_Sorter100|10273_ , \new_Sorter100|10274_ ,
    \new_Sorter100|10275_ , \new_Sorter100|10276_ , \new_Sorter100|10277_ ,
    \new_Sorter100|10278_ , \new_Sorter100|10279_ , \new_Sorter100|10280_ ,
    \new_Sorter100|10281_ , \new_Sorter100|10282_ , \new_Sorter100|10283_ ,
    \new_Sorter100|10284_ , \new_Sorter100|10285_ , \new_Sorter100|10286_ ,
    \new_Sorter100|10287_ , \new_Sorter100|10288_ , \new_Sorter100|10289_ ,
    \new_Sorter100|10290_ , \new_Sorter100|10291_ , \new_Sorter100|10292_ ,
    \new_Sorter100|10293_ , \new_Sorter100|10294_ , \new_Sorter100|10295_ ,
    \new_Sorter100|10296_ , \new_Sorter100|10297_ , \new_Sorter100|10298_ ,
    \new_Sorter100|10299_ , \new_Sorter100|10300_ , \new_Sorter100|10399_ ,
    \new_Sorter100|10301_ , \new_Sorter100|10302_ , \new_Sorter100|10303_ ,
    \new_Sorter100|10304_ , \new_Sorter100|10305_ , \new_Sorter100|10306_ ,
    \new_Sorter100|10307_ , \new_Sorter100|10308_ , \new_Sorter100|10309_ ,
    \new_Sorter100|10310_ , \new_Sorter100|10311_ , \new_Sorter100|10312_ ,
    \new_Sorter100|10313_ , \new_Sorter100|10314_ , \new_Sorter100|10315_ ,
    \new_Sorter100|10316_ , \new_Sorter100|10317_ , \new_Sorter100|10318_ ,
    \new_Sorter100|10319_ , \new_Sorter100|10320_ , \new_Sorter100|10321_ ,
    \new_Sorter100|10322_ , \new_Sorter100|10323_ , \new_Sorter100|10324_ ,
    \new_Sorter100|10325_ , \new_Sorter100|10326_ , \new_Sorter100|10327_ ,
    \new_Sorter100|10328_ , \new_Sorter100|10329_ , \new_Sorter100|10330_ ,
    \new_Sorter100|10331_ , \new_Sorter100|10332_ , \new_Sorter100|10333_ ,
    \new_Sorter100|10334_ , \new_Sorter100|10335_ , \new_Sorter100|10336_ ,
    \new_Sorter100|10337_ , \new_Sorter100|10338_ , \new_Sorter100|10339_ ,
    \new_Sorter100|10340_ , \new_Sorter100|10341_ , \new_Sorter100|10342_ ,
    \new_Sorter100|10343_ , \new_Sorter100|10344_ , \new_Sorter100|10345_ ,
    \new_Sorter100|10346_ , \new_Sorter100|10347_ , \new_Sorter100|10348_ ,
    \new_Sorter100|10349_ , \new_Sorter100|10350_ , \new_Sorter100|10351_ ,
    \new_Sorter100|10352_ , \new_Sorter100|10353_ , \new_Sorter100|10354_ ,
    \new_Sorter100|10355_ , \new_Sorter100|10356_ , \new_Sorter100|10357_ ,
    \new_Sorter100|10358_ , \new_Sorter100|10359_ , \new_Sorter100|10360_ ,
    \new_Sorter100|10361_ , \new_Sorter100|10362_ , \new_Sorter100|10363_ ,
    \new_Sorter100|10364_ , \new_Sorter100|10365_ , \new_Sorter100|10366_ ,
    \new_Sorter100|10367_ , \new_Sorter100|10368_ , \new_Sorter100|10369_ ,
    \new_Sorter100|10370_ , \new_Sorter100|10371_ , \new_Sorter100|10372_ ,
    \new_Sorter100|10373_ , \new_Sorter100|10374_ , \new_Sorter100|10375_ ,
    \new_Sorter100|10376_ , \new_Sorter100|10377_ , \new_Sorter100|10378_ ,
    \new_Sorter100|10379_ , \new_Sorter100|10380_ , \new_Sorter100|10381_ ,
    \new_Sorter100|10382_ , \new_Sorter100|10383_ , \new_Sorter100|10384_ ,
    \new_Sorter100|10385_ , \new_Sorter100|10386_ , \new_Sorter100|10387_ ,
    \new_Sorter100|10388_ , \new_Sorter100|10389_ , \new_Sorter100|10390_ ,
    \new_Sorter100|10391_ , \new_Sorter100|10392_ , \new_Sorter100|10393_ ,
    \new_Sorter100|10394_ , \new_Sorter100|10395_ , \new_Sorter100|10396_ ,
    \new_Sorter100|10397_ , \new_Sorter100|10398_ , \new_Sorter100|10400_ ,
    \new_Sorter100|10401_ , \new_Sorter100|10402_ , \new_Sorter100|10403_ ,
    \new_Sorter100|10404_ , \new_Sorter100|10405_ , \new_Sorter100|10406_ ,
    \new_Sorter100|10407_ , \new_Sorter100|10408_ , \new_Sorter100|10409_ ,
    \new_Sorter100|10410_ , \new_Sorter100|10411_ , \new_Sorter100|10412_ ,
    \new_Sorter100|10413_ , \new_Sorter100|10414_ , \new_Sorter100|10415_ ,
    \new_Sorter100|10416_ , \new_Sorter100|10417_ , \new_Sorter100|10418_ ,
    \new_Sorter100|10419_ , \new_Sorter100|10420_ , \new_Sorter100|10421_ ,
    \new_Sorter100|10422_ , \new_Sorter100|10423_ , \new_Sorter100|10424_ ,
    \new_Sorter100|10425_ , \new_Sorter100|10426_ , \new_Sorter100|10427_ ,
    \new_Sorter100|10428_ , \new_Sorter100|10429_ , \new_Sorter100|10430_ ,
    \new_Sorter100|10431_ , \new_Sorter100|10432_ , \new_Sorter100|10433_ ,
    \new_Sorter100|10434_ , \new_Sorter100|10435_ , \new_Sorter100|10436_ ,
    \new_Sorter100|10437_ , \new_Sorter100|10438_ , \new_Sorter100|10439_ ,
    \new_Sorter100|10440_ , \new_Sorter100|10441_ , \new_Sorter100|10442_ ,
    \new_Sorter100|10443_ , \new_Sorter100|10444_ , \new_Sorter100|10445_ ,
    \new_Sorter100|10446_ , \new_Sorter100|10447_ , \new_Sorter100|10448_ ,
    \new_Sorter100|10449_ , \new_Sorter100|10450_ , \new_Sorter100|10451_ ,
    \new_Sorter100|10452_ , \new_Sorter100|10453_ , \new_Sorter100|10454_ ,
    \new_Sorter100|10455_ , \new_Sorter100|10456_ , \new_Sorter100|10457_ ,
    \new_Sorter100|10458_ , \new_Sorter100|10459_ , \new_Sorter100|10460_ ,
    \new_Sorter100|10461_ , \new_Sorter100|10462_ , \new_Sorter100|10463_ ,
    \new_Sorter100|10464_ , \new_Sorter100|10465_ , \new_Sorter100|10466_ ,
    \new_Sorter100|10467_ , \new_Sorter100|10468_ , \new_Sorter100|10469_ ,
    \new_Sorter100|10470_ , \new_Sorter100|10471_ , \new_Sorter100|10472_ ,
    \new_Sorter100|10473_ , \new_Sorter100|10474_ , \new_Sorter100|10475_ ,
    \new_Sorter100|10476_ , \new_Sorter100|10477_ , \new_Sorter100|10478_ ,
    \new_Sorter100|10479_ , \new_Sorter100|10480_ , \new_Sorter100|10481_ ,
    \new_Sorter100|10482_ , \new_Sorter100|10483_ , \new_Sorter100|10484_ ,
    \new_Sorter100|10485_ , \new_Sorter100|10486_ , \new_Sorter100|10487_ ,
    \new_Sorter100|10488_ , \new_Sorter100|10489_ , \new_Sorter100|10490_ ,
    \new_Sorter100|10491_ , \new_Sorter100|10492_ , \new_Sorter100|10493_ ,
    \new_Sorter100|10494_ , \new_Sorter100|10495_ , \new_Sorter100|10496_ ,
    \new_Sorter100|10497_ , \new_Sorter100|10498_ , \new_Sorter100|10499_ ,
    \new_Sorter100|10500_ , \new_Sorter100|10599_ , \new_Sorter100|10501_ ,
    \new_Sorter100|10502_ , \new_Sorter100|10503_ , \new_Sorter100|10504_ ,
    \new_Sorter100|10505_ , \new_Sorter100|10506_ , \new_Sorter100|10507_ ,
    \new_Sorter100|10508_ , \new_Sorter100|10509_ , \new_Sorter100|10510_ ,
    \new_Sorter100|10511_ , \new_Sorter100|10512_ , \new_Sorter100|10513_ ,
    \new_Sorter100|10514_ , \new_Sorter100|10515_ , \new_Sorter100|10516_ ,
    \new_Sorter100|10517_ , \new_Sorter100|10518_ , \new_Sorter100|10519_ ,
    \new_Sorter100|10520_ , \new_Sorter100|10521_ , \new_Sorter100|10522_ ,
    \new_Sorter100|10523_ , \new_Sorter100|10524_ , \new_Sorter100|10525_ ,
    \new_Sorter100|10526_ , \new_Sorter100|10527_ , \new_Sorter100|10528_ ,
    \new_Sorter100|10529_ , \new_Sorter100|10530_ , \new_Sorter100|10531_ ,
    \new_Sorter100|10532_ , \new_Sorter100|10533_ , \new_Sorter100|10534_ ,
    \new_Sorter100|10535_ , \new_Sorter100|10536_ , \new_Sorter100|10537_ ,
    \new_Sorter100|10538_ , \new_Sorter100|10539_ , \new_Sorter100|10540_ ,
    \new_Sorter100|10541_ , \new_Sorter100|10542_ , \new_Sorter100|10543_ ,
    \new_Sorter100|10544_ , \new_Sorter100|10545_ , \new_Sorter100|10546_ ,
    \new_Sorter100|10547_ , \new_Sorter100|10548_ , \new_Sorter100|10549_ ,
    \new_Sorter100|10550_ , \new_Sorter100|10551_ , \new_Sorter100|10552_ ,
    \new_Sorter100|10553_ , \new_Sorter100|10554_ , \new_Sorter100|10555_ ,
    \new_Sorter100|10556_ , \new_Sorter100|10557_ , \new_Sorter100|10558_ ,
    \new_Sorter100|10559_ , \new_Sorter100|10560_ , \new_Sorter100|10561_ ,
    \new_Sorter100|10562_ , \new_Sorter100|10563_ , \new_Sorter100|10564_ ,
    \new_Sorter100|10565_ , \new_Sorter100|10566_ , \new_Sorter100|10567_ ,
    \new_Sorter100|10568_ , \new_Sorter100|10569_ , \new_Sorter100|10570_ ,
    \new_Sorter100|10571_ , \new_Sorter100|10572_ , \new_Sorter100|10573_ ,
    \new_Sorter100|10574_ , \new_Sorter100|10575_ , \new_Sorter100|10576_ ,
    \new_Sorter100|10577_ , \new_Sorter100|10578_ , \new_Sorter100|10579_ ,
    \new_Sorter100|10580_ , \new_Sorter100|10581_ , \new_Sorter100|10582_ ,
    \new_Sorter100|10583_ , \new_Sorter100|10584_ , \new_Sorter100|10585_ ,
    \new_Sorter100|10586_ , \new_Sorter100|10587_ , \new_Sorter100|10588_ ,
    \new_Sorter100|10589_ , \new_Sorter100|10590_ , \new_Sorter100|10591_ ,
    \new_Sorter100|10592_ , \new_Sorter100|10593_ , \new_Sorter100|10594_ ,
    \new_Sorter100|10595_ , \new_Sorter100|10596_ , \new_Sorter100|10597_ ,
    \new_Sorter100|10598_ , \new_Sorter100|10600_ , \new_Sorter100|10601_ ,
    \new_Sorter100|10602_ , \new_Sorter100|10603_ , \new_Sorter100|10604_ ,
    \new_Sorter100|10605_ , \new_Sorter100|10606_ , \new_Sorter100|10607_ ,
    \new_Sorter100|10608_ , \new_Sorter100|10609_ , \new_Sorter100|10610_ ,
    \new_Sorter100|10611_ , \new_Sorter100|10612_ , \new_Sorter100|10613_ ,
    \new_Sorter100|10614_ , \new_Sorter100|10615_ , \new_Sorter100|10616_ ,
    \new_Sorter100|10617_ , \new_Sorter100|10618_ , \new_Sorter100|10619_ ,
    \new_Sorter100|10620_ , \new_Sorter100|10621_ , \new_Sorter100|10622_ ,
    \new_Sorter100|10623_ , \new_Sorter100|10624_ , \new_Sorter100|10625_ ,
    \new_Sorter100|10626_ , \new_Sorter100|10627_ , \new_Sorter100|10628_ ,
    \new_Sorter100|10629_ , \new_Sorter100|10630_ , \new_Sorter100|10631_ ,
    \new_Sorter100|10632_ , \new_Sorter100|10633_ , \new_Sorter100|10634_ ,
    \new_Sorter100|10635_ , \new_Sorter100|10636_ , \new_Sorter100|10637_ ,
    \new_Sorter100|10638_ , \new_Sorter100|10639_ , \new_Sorter100|10640_ ,
    \new_Sorter100|10641_ , \new_Sorter100|10642_ , \new_Sorter100|10643_ ,
    \new_Sorter100|10644_ , \new_Sorter100|10645_ , \new_Sorter100|10646_ ,
    \new_Sorter100|10647_ , \new_Sorter100|10648_ , \new_Sorter100|10649_ ,
    \new_Sorter100|10650_ , \new_Sorter100|10651_ , \new_Sorter100|10652_ ,
    \new_Sorter100|10653_ , \new_Sorter100|10654_ , \new_Sorter100|10655_ ,
    \new_Sorter100|10656_ , \new_Sorter100|10657_ , \new_Sorter100|10658_ ,
    \new_Sorter100|10659_ , \new_Sorter100|10660_ , \new_Sorter100|10661_ ,
    \new_Sorter100|10662_ , \new_Sorter100|10663_ , \new_Sorter100|10664_ ,
    \new_Sorter100|10665_ , \new_Sorter100|10666_ , \new_Sorter100|10667_ ,
    \new_Sorter100|10668_ , \new_Sorter100|10669_ , \new_Sorter100|10670_ ,
    \new_Sorter100|10671_ , \new_Sorter100|10672_ , \new_Sorter100|10673_ ,
    \new_Sorter100|10674_ , \new_Sorter100|10675_ , \new_Sorter100|10676_ ,
    \new_Sorter100|10677_ , \new_Sorter100|10678_ , \new_Sorter100|10679_ ,
    \new_Sorter100|10680_ , \new_Sorter100|10681_ , \new_Sorter100|10682_ ,
    \new_Sorter100|10683_ , \new_Sorter100|10684_ , \new_Sorter100|10685_ ,
    \new_Sorter100|10686_ , \new_Sorter100|10687_ , \new_Sorter100|10688_ ,
    \new_Sorter100|10689_ , \new_Sorter100|10690_ , \new_Sorter100|10691_ ,
    \new_Sorter100|10692_ , \new_Sorter100|10693_ , \new_Sorter100|10694_ ,
    \new_Sorter100|10695_ , \new_Sorter100|10696_ , \new_Sorter100|10697_ ,
    \new_Sorter100|10698_ , \new_Sorter100|10699_ , \new_Sorter100|10700_ ,
    \new_Sorter100|10799_ , \new_Sorter100|10701_ , \new_Sorter100|10702_ ,
    \new_Sorter100|10703_ , \new_Sorter100|10704_ , \new_Sorter100|10705_ ,
    \new_Sorter100|10706_ , \new_Sorter100|10707_ , \new_Sorter100|10708_ ,
    \new_Sorter100|10709_ , \new_Sorter100|10710_ , \new_Sorter100|10711_ ,
    \new_Sorter100|10712_ , \new_Sorter100|10713_ , \new_Sorter100|10714_ ,
    \new_Sorter100|10715_ , \new_Sorter100|10716_ , \new_Sorter100|10717_ ,
    \new_Sorter100|10718_ , \new_Sorter100|10719_ , \new_Sorter100|10720_ ,
    \new_Sorter100|10721_ , \new_Sorter100|10722_ , \new_Sorter100|10723_ ,
    \new_Sorter100|10724_ , \new_Sorter100|10725_ , \new_Sorter100|10726_ ,
    \new_Sorter100|10727_ , \new_Sorter100|10728_ , \new_Sorter100|10729_ ,
    \new_Sorter100|10730_ , \new_Sorter100|10731_ , \new_Sorter100|10732_ ,
    \new_Sorter100|10733_ , \new_Sorter100|10734_ , \new_Sorter100|10735_ ,
    \new_Sorter100|10736_ , \new_Sorter100|10737_ , \new_Sorter100|10738_ ,
    \new_Sorter100|10739_ , \new_Sorter100|10740_ , \new_Sorter100|10741_ ,
    \new_Sorter100|10742_ , \new_Sorter100|10743_ , \new_Sorter100|10744_ ,
    \new_Sorter100|10745_ , \new_Sorter100|10746_ , \new_Sorter100|10747_ ,
    \new_Sorter100|10748_ , \new_Sorter100|10749_ , \new_Sorter100|10750_ ,
    \new_Sorter100|10751_ , \new_Sorter100|10752_ , \new_Sorter100|10753_ ,
    \new_Sorter100|10754_ , \new_Sorter100|10755_ , \new_Sorter100|10756_ ,
    \new_Sorter100|10757_ , \new_Sorter100|10758_ , \new_Sorter100|10759_ ,
    \new_Sorter100|10760_ , \new_Sorter100|10761_ , \new_Sorter100|10762_ ,
    \new_Sorter100|10763_ , \new_Sorter100|10764_ , \new_Sorter100|10765_ ,
    \new_Sorter100|10766_ , \new_Sorter100|10767_ , \new_Sorter100|10768_ ,
    \new_Sorter100|10769_ , \new_Sorter100|10770_ , \new_Sorter100|10771_ ,
    \new_Sorter100|10772_ , \new_Sorter100|10773_ , \new_Sorter100|10774_ ,
    \new_Sorter100|10775_ , \new_Sorter100|10776_ , \new_Sorter100|10777_ ,
    \new_Sorter100|10778_ , \new_Sorter100|10779_ , \new_Sorter100|10780_ ,
    \new_Sorter100|10781_ , \new_Sorter100|10782_ , \new_Sorter100|10783_ ,
    \new_Sorter100|10784_ , \new_Sorter100|10785_ , \new_Sorter100|10786_ ,
    \new_Sorter100|10787_ , \new_Sorter100|10788_ , \new_Sorter100|10789_ ,
    \new_Sorter100|10790_ , \new_Sorter100|10791_ , \new_Sorter100|10792_ ,
    \new_Sorter100|10793_ , \new_Sorter100|10794_ , \new_Sorter100|10795_ ,
    \new_Sorter100|10796_ , \new_Sorter100|10797_ , \new_Sorter100|10798_ ,
    \new_Sorter100|10800_ , \new_Sorter100|10801_ , \new_Sorter100|10802_ ,
    \new_Sorter100|10803_ , \new_Sorter100|10804_ , \new_Sorter100|10805_ ,
    \new_Sorter100|10806_ , \new_Sorter100|10807_ , \new_Sorter100|10808_ ,
    \new_Sorter100|10809_ , \new_Sorter100|10810_ , \new_Sorter100|10811_ ,
    \new_Sorter100|10812_ , \new_Sorter100|10813_ , \new_Sorter100|10814_ ,
    \new_Sorter100|10815_ , \new_Sorter100|10816_ , \new_Sorter100|10817_ ,
    \new_Sorter100|10818_ , \new_Sorter100|10819_ , \new_Sorter100|10820_ ,
    \new_Sorter100|10821_ , \new_Sorter100|10822_ , \new_Sorter100|10823_ ,
    \new_Sorter100|10824_ , \new_Sorter100|10825_ , \new_Sorter100|10826_ ,
    \new_Sorter100|10827_ , \new_Sorter100|10828_ , \new_Sorter100|10829_ ,
    \new_Sorter100|10830_ , \new_Sorter100|10831_ , \new_Sorter100|10832_ ,
    \new_Sorter100|10833_ , \new_Sorter100|10834_ , \new_Sorter100|10835_ ,
    \new_Sorter100|10836_ , \new_Sorter100|10837_ , \new_Sorter100|10838_ ,
    \new_Sorter100|10839_ , \new_Sorter100|10840_ , \new_Sorter100|10841_ ,
    \new_Sorter100|10842_ , \new_Sorter100|10843_ , \new_Sorter100|10844_ ,
    \new_Sorter100|10845_ , \new_Sorter100|10846_ , \new_Sorter100|10847_ ,
    \new_Sorter100|10848_ , \new_Sorter100|10849_ , \new_Sorter100|10850_ ,
    \new_Sorter100|10851_ , \new_Sorter100|10852_ , \new_Sorter100|10853_ ,
    \new_Sorter100|10854_ , \new_Sorter100|10855_ , \new_Sorter100|10856_ ,
    \new_Sorter100|10857_ , \new_Sorter100|10858_ , \new_Sorter100|10859_ ,
    \new_Sorter100|10860_ , \new_Sorter100|10861_ , \new_Sorter100|10862_ ,
    \new_Sorter100|10863_ , \new_Sorter100|10864_ , \new_Sorter100|10865_ ,
    \new_Sorter100|10866_ , \new_Sorter100|10867_ , \new_Sorter100|10868_ ,
    \new_Sorter100|10869_ , \new_Sorter100|10870_ , \new_Sorter100|10871_ ,
    \new_Sorter100|10872_ , \new_Sorter100|10873_ , \new_Sorter100|10874_ ,
    \new_Sorter100|10875_ , \new_Sorter100|10876_ , \new_Sorter100|10877_ ,
    \new_Sorter100|10878_ , \new_Sorter100|10879_ , \new_Sorter100|10880_ ,
    \new_Sorter100|10881_ , \new_Sorter100|10882_ , \new_Sorter100|10883_ ,
    \new_Sorter100|10884_ , \new_Sorter100|10885_ , \new_Sorter100|10886_ ,
    \new_Sorter100|10887_ , \new_Sorter100|10888_ , \new_Sorter100|10889_ ,
    \new_Sorter100|10890_ , \new_Sorter100|10891_ , \new_Sorter100|10892_ ,
    \new_Sorter100|10893_ , \new_Sorter100|10894_ , \new_Sorter100|10895_ ,
    \new_Sorter100|10896_ , \new_Sorter100|10897_ , \new_Sorter100|10898_ ,
    \new_Sorter100|10899_ , \new_Sorter100|10900_ , \new_Sorter100|10999_ ,
    \new_Sorter100|10901_ , \new_Sorter100|10902_ , \new_Sorter100|10903_ ,
    \new_Sorter100|10904_ , \new_Sorter100|10905_ , \new_Sorter100|10906_ ,
    \new_Sorter100|10907_ , \new_Sorter100|10908_ , \new_Sorter100|10909_ ,
    \new_Sorter100|10910_ , \new_Sorter100|10911_ , \new_Sorter100|10912_ ,
    \new_Sorter100|10913_ , \new_Sorter100|10914_ , \new_Sorter100|10915_ ,
    \new_Sorter100|10916_ , \new_Sorter100|10917_ , \new_Sorter100|10918_ ,
    \new_Sorter100|10919_ , \new_Sorter100|10920_ , \new_Sorter100|10921_ ,
    \new_Sorter100|10922_ , \new_Sorter100|10923_ , \new_Sorter100|10924_ ,
    \new_Sorter100|10925_ , \new_Sorter100|10926_ , \new_Sorter100|10927_ ,
    \new_Sorter100|10928_ , \new_Sorter100|10929_ , \new_Sorter100|10930_ ,
    \new_Sorter100|10931_ , \new_Sorter100|10932_ , \new_Sorter100|10933_ ,
    \new_Sorter100|10934_ , \new_Sorter100|10935_ , \new_Sorter100|10936_ ,
    \new_Sorter100|10937_ , \new_Sorter100|10938_ , \new_Sorter100|10939_ ,
    \new_Sorter100|10940_ , \new_Sorter100|10941_ , \new_Sorter100|10942_ ,
    \new_Sorter100|10943_ , \new_Sorter100|10944_ , \new_Sorter100|10945_ ,
    \new_Sorter100|10946_ , \new_Sorter100|10947_ , \new_Sorter100|10948_ ,
    \new_Sorter100|10949_ , \new_Sorter100|10950_ , \new_Sorter100|10951_ ,
    \new_Sorter100|10952_ , \new_Sorter100|10953_ , \new_Sorter100|10954_ ,
    \new_Sorter100|10955_ , \new_Sorter100|10956_ , \new_Sorter100|10957_ ,
    \new_Sorter100|10958_ , \new_Sorter100|10959_ , \new_Sorter100|10960_ ,
    \new_Sorter100|10961_ , \new_Sorter100|10962_ , \new_Sorter100|10963_ ,
    \new_Sorter100|10964_ , \new_Sorter100|10965_ , \new_Sorter100|10966_ ,
    \new_Sorter100|10967_ , \new_Sorter100|10968_ , \new_Sorter100|10969_ ,
    \new_Sorter100|10970_ , \new_Sorter100|10971_ , \new_Sorter100|10972_ ,
    \new_Sorter100|10973_ , \new_Sorter100|10974_ , \new_Sorter100|10975_ ,
    \new_Sorter100|10976_ , \new_Sorter100|10977_ , \new_Sorter100|10978_ ,
    \new_Sorter100|10979_ , \new_Sorter100|10980_ , \new_Sorter100|10981_ ,
    \new_Sorter100|10982_ , \new_Sorter100|10983_ , \new_Sorter100|10984_ ,
    \new_Sorter100|10985_ , \new_Sorter100|10986_ , \new_Sorter100|10987_ ,
    \new_Sorter100|10988_ , \new_Sorter100|10989_ , \new_Sorter100|10990_ ,
    \new_Sorter100|10991_ , \new_Sorter100|10992_ , \new_Sorter100|10993_ ,
    \new_Sorter100|10994_ , \new_Sorter100|10995_ , \new_Sorter100|10996_ ,
    \new_Sorter100|10997_ , \new_Sorter100|10998_ , \new_Sorter100|11000_ ,
    \new_Sorter100|11001_ , \new_Sorter100|11002_ , \new_Sorter100|11003_ ,
    \new_Sorter100|11004_ , \new_Sorter100|11005_ , \new_Sorter100|11006_ ,
    \new_Sorter100|11007_ , \new_Sorter100|11008_ , \new_Sorter100|11009_ ,
    \new_Sorter100|11010_ , \new_Sorter100|11011_ , \new_Sorter100|11012_ ,
    \new_Sorter100|11013_ , \new_Sorter100|11014_ , \new_Sorter100|11015_ ,
    \new_Sorter100|11016_ , \new_Sorter100|11017_ , \new_Sorter100|11018_ ,
    \new_Sorter100|11019_ , \new_Sorter100|11020_ , \new_Sorter100|11021_ ,
    \new_Sorter100|11022_ , \new_Sorter100|11023_ , \new_Sorter100|11024_ ,
    \new_Sorter100|11025_ , \new_Sorter100|11026_ , \new_Sorter100|11027_ ,
    \new_Sorter100|11028_ , \new_Sorter100|11029_ , \new_Sorter100|11030_ ,
    \new_Sorter100|11031_ , \new_Sorter100|11032_ , \new_Sorter100|11033_ ,
    \new_Sorter100|11034_ , \new_Sorter100|11035_ , \new_Sorter100|11036_ ,
    \new_Sorter100|11037_ , \new_Sorter100|11038_ , \new_Sorter100|11039_ ,
    \new_Sorter100|11040_ , \new_Sorter100|11041_ , \new_Sorter100|11042_ ,
    \new_Sorter100|11043_ , \new_Sorter100|11044_ , \new_Sorter100|11045_ ,
    \new_Sorter100|11046_ , \new_Sorter100|11047_ , \new_Sorter100|11048_ ,
    \new_Sorter100|11049_ , \new_Sorter100|11050_ , \new_Sorter100|11051_ ,
    \new_Sorter100|11052_ , \new_Sorter100|11053_ , \new_Sorter100|11054_ ,
    \new_Sorter100|11055_ , \new_Sorter100|11056_ , \new_Sorter100|11057_ ,
    \new_Sorter100|11058_ , \new_Sorter100|11059_ , \new_Sorter100|11060_ ,
    \new_Sorter100|11061_ , \new_Sorter100|11062_ , \new_Sorter100|11063_ ,
    \new_Sorter100|11064_ , \new_Sorter100|11065_ , \new_Sorter100|11066_ ,
    \new_Sorter100|11067_ , \new_Sorter100|11068_ , \new_Sorter100|11069_ ,
    \new_Sorter100|11070_ , \new_Sorter100|11071_ , \new_Sorter100|11072_ ,
    \new_Sorter100|11073_ , \new_Sorter100|11074_ , \new_Sorter100|11075_ ,
    \new_Sorter100|11076_ , \new_Sorter100|11077_ , \new_Sorter100|11078_ ,
    \new_Sorter100|11079_ , \new_Sorter100|11080_ , \new_Sorter100|11081_ ,
    \new_Sorter100|11082_ , \new_Sorter100|11083_ , \new_Sorter100|11084_ ,
    \new_Sorter100|11085_ , \new_Sorter100|11086_ , \new_Sorter100|11087_ ,
    \new_Sorter100|11088_ , \new_Sorter100|11089_ , \new_Sorter100|11090_ ,
    \new_Sorter100|11091_ , \new_Sorter100|11092_ , \new_Sorter100|11093_ ,
    \new_Sorter100|11094_ , \new_Sorter100|11095_ , \new_Sorter100|11096_ ,
    \new_Sorter100|11097_ , \new_Sorter100|11098_ , \new_Sorter100|11099_ ,
    \new_Sorter100|11100_ , \new_Sorter100|11199_ , \new_Sorter100|11101_ ,
    \new_Sorter100|11102_ , \new_Sorter100|11103_ , \new_Sorter100|11104_ ,
    \new_Sorter100|11105_ , \new_Sorter100|11106_ , \new_Sorter100|11107_ ,
    \new_Sorter100|11108_ , \new_Sorter100|11109_ , \new_Sorter100|11110_ ,
    \new_Sorter100|11111_ , \new_Sorter100|11112_ , \new_Sorter100|11113_ ,
    \new_Sorter100|11114_ , \new_Sorter100|11115_ , \new_Sorter100|11116_ ,
    \new_Sorter100|11117_ , \new_Sorter100|11118_ , \new_Sorter100|11119_ ,
    \new_Sorter100|11120_ , \new_Sorter100|11121_ , \new_Sorter100|11122_ ,
    \new_Sorter100|11123_ , \new_Sorter100|11124_ , \new_Sorter100|11125_ ,
    \new_Sorter100|11126_ , \new_Sorter100|11127_ , \new_Sorter100|11128_ ,
    \new_Sorter100|11129_ , \new_Sorter100|11130_ , \new_Sorter100|11131_ ,
    \new_Sorter100|11132_ , \new_Sorter100|11133_ , \new_Sorter100|11134_ ,
    \new_Sorter100|11135_ , \new_Sorter100|11136_ , \new_Sorter100|11137_ ,
    \new_Sorter100|11138_ , \new_Sorter100|11139_ , \new_Sorter100|11140_ ,
    \new_Sorter100|11141_ , \new_Sorter100|11142_ , \new_Sorter100|11143_ ,
    \new_Sorter100|11144_ , \new_Sorter100|11145_ , \new_Sorter100|11146_ ,
    \new_Sorter100|11147_ , \new_Sorter100|11148_ , \new_Sorter100|11149_ ,
    \new_Sorter100|11150_ , \new_Sorter100|11151_ , \new_Sorter100|11152_ ,
    \new_Sorter100|11153_ , \new_Sorter100|11154_ , \new_Sorter100|11155_ ,
    \new_Sorter100|11156_ , \new_Sorter100|11157_ , \new_Sorter100|11158_ ,
    \new_Sorter100|11159_ , \new_Sorter100|11160_ , \new_Sorter100|11161_ ,
    \new_Sorter100|11162_ , \new_Sorter100|11163_ , \new_Sorter100|11164_ ,
    \new_Sorter100|11165_ , \new_Sorter100|11166_ , \new_Sorter100|11167_ ,
    \new_Sorter100|11168_ , \new_Sorter100|11169_ , \new_Sorter100|11170_ ,
    \new_Sorter100|11171_ , \new_Sorter100|11172_ , \new_Sorter100|11173_ ,
    \new_Sorter100|11174_ , \new_Sorter100|11175_ , \new_Sorter100|11176_ ,
    \new_Sorter100|11177_ , \new_Sorter100|11178_ , \new_Sorter100|11179_ ,
    \new_Sorter100|11180_ , \new_Sorter100|11181_ , \new_Sorter100|11182_ ,
    \new_Sorter100|11183_ , \new_Sorter100|11184_ , \new_Sorter100|11185_ ,
    \new_Sorter100|11186_ , \new_Sorter100|11187_ , \new_Sorter100|11188_ ,
    \new_Sorter100|11189_ , \new_Sorter100|11190_ , \new_Sorter100|11191_ ,
    \new_Sorter100|11192_ , \new_Sorter100|11193_ , \new_Sorter100|11194_ ,
    \new_Sorter100|11195_ , \new_Sorter100|11196_ , \new_Sorter100|11197_ ,
    \new_Sorter100|11198_ , \new_Sorter100|11200_ , \new_Sorter100|11201_ ,
    \new_Sorter100|11202_ , \new_Sorter100|11203_ , \new_Sorter100|11204_ ,
    \new_Sorter100|11205_ , \new_Sorter100|11206_ , \new_Sorter100|11207_ ,
    \new_Sorter100|11208_ , \new_Sorter100|11209_ , \new_Sorter100|11210_ ,
    \new_Sorter100|11211_ , \new_Sorter100|11212_ , \new_Sorter100|11213_ ,
    \new_Sorter100|11214_ , \new_Sorter100|11215_ , \new_Sorter100|11216_ ,
    \new_Sorter100|11217_ , \new_Sorter100|11218_ , \new_Sorter100|11219_ ,
    \new_Sorter100|11220_ , \new_Sorter100|11221_ , \new_Sorter100|11222_ ,
    \new_Sorter100|11223_ , \new_Sorter100|11224_ , \new_Sorter100|11225_ ,
    \new_Sorter100|11226_ , \new_Sorter100|11227_ , \new_Sorter100|11228_ ,
    \new_Sorter100|11229_ , \new_Sorter100|11230_ , \new_Sorter100|11231_ ,
    \new_Sorter100|11232_ , \new_Sorter100|11233_ , \new_Sorter100|11234_ ,
    \new_Sorter100|11235_ , \new_Sorter100|11236_ , \new_Sorter100|11237_ ,
    \new_Sorter100|11238_ , \new_Sorter100|11239_ , \new_Sorter100|11240_ ,
    \new_Sorter100|11241_ , \new_Sorter100|11242_ , \new_Sorter100|11243_ ,
    \new_Sorter100|11244_ , \new_Sorter100|11245_ , \new_Sorter100|11246_ ,
    \new_Sorter100|11247_ , \new_Sorter100|11248_ , \new_Sorter100|11249_ ,
    \new_Sorter100|11250_ , \new_Sorter100|11251_ , \new_Sorter100|11252_ ,
    \new_Sorter100|11253_ , \new_Sorter100|11254_ , \new_Sorter100|11255_ ,
    \new_Sorter100|11256_ , \new_Sorter100|11257_ , \new_Sorter100|11258_ ,
    \new_Sorter100|11259_ , \new_Sorter100|11260_ , \new_Sorter100|11261_ ,
    \new_Sorter100|11262_ , \new_Sorter100|11263_ , \new_Sorter100|11264_ ,
    \new_Sorter100|11265_ , \new_Sorter100|11266_ , \new_Sorter100|11267_ ,
    \new_Sorter100|11268_ , \new_Sorter100|11269_ , \new_Sorter100|11270_ ,
    \new_Sorter100|11271_ , \new_Sorter100|11272_ , \new_Sorter100|11273_ ,
    \new_Sorter100|11274_ , \new_Sorter100|11275_ , \new_Sorter100|11276_ ,
    \new_Sorter100|11277_ , \new_Sorter100|11278_ , \new_Sorter100|11279_ ,
    \new_Sorter100|11280_ , \new_Sorter100|11281_ , \new_Sorter100|11282_ ,
    \new_Sorter100|11283_ , \new_Sorter100|11284_ , \new_Sorter100|11285_ ,
    \new_Sorter100|11286_ , \new_Sorter100|11287_ , \new_Sorter100|11288_ ,
    \new_Sorter100|11289_ , \new_Sorter100|11290_ , \new_Sorter100|11291_ ,
    \new_Sorter100|11292_ , \new_Sorter100|11293_ , \new_Sorter100|11294_ ,
    \new_Sorter100|11295_ , \new_Sorter100|11296_ , \new_Sorter100|11297_ ,
    \new_Sorter100|11298_ , \new_Sorter100|11299_ , \new_Sorter100|11300_ ,
    \new_Sorter100|11399_ , \new_Sorter100|11301_ , \new_Sorter100|11302_ ,
    \new_Sorter100|11303_ , \new_Sorter100|11304_ , \new_Sorter100|11305_ ,
    \new_Sorter100|11306_ , \new_Sorter100|11307_ , \new_Sorter100|11308_ ,
    \new_Sorter100|11309_ , \new_Sorter100|11310_ , \new_Sorter100|11311_ ,
    \new_Sorter100|11312_ , \new_Sorter100|11313_ , \new_Sorter100|11314_ ,
    \new_Sorter100|11315_ , \new_Sorter100|11316_ , \new_Sorter100|11317_ ,
    \new_Sorter100|11318_ , \new_Sorter100|11319_ , \new_Sorter100|11320_ ,
    \new_Sorter100|11321_ , \new_Sorter100|11322_ , \new_Sorter100|11323_ ,
    \new_Sorter100|11324_ , \new_Sorter100|11325_ , \new_Sorter100|11326_ ,
    \new_Sorter100|11327_ , \new_Sorter100|11328_ , \new_Sorter100|11329_ ,
    \new_Sorter100|11330_ , \new_Sorter100|11331_ , \new_Sorter100|11332_ ,
    \new_Sorter100|11333_ , \new_Sorter100|11334_ , \new_Sorter100|11335_ ,
    \new_Sorter100|11336_ , \new_Sorter100|11337_ , \new_Sorter100|11338_ ,
    \new_Sorter100|11339_ , \new_Sorter100|11340_ , \new_Sorter100|11341_ ,
    \new_Sorter100|11342_ , \new_Sorter100|11343_ , \new_Sorter100|11344_ ,
    \new_Sorter100|11345_ , \new_Sorter100|11346_ , \new_Sorter100|11347_ ,
    \new_Sorter100|11348_ , \new_Sorter100|11349_ , \new_Sorter100|11350_ ,
    \new_Sorter100|11351_ , \new_Sorter100|11352_ , \new_Sorter100|11353_ ,
    \new_Sorter100|11354_ , \new_Sorter100|11355_ , \new_Sorter100|11356_ ,
    \new_Sorter100|11357_ , \new_Sorter100|11358_ , \new_Sorter100|11359_ ,
    \new_Sorter100|11360_ , \new_Sorter100|11361_ , \new_Sorter100|11362_ ,
    \new_Sorter100|11363_ , \new_Sorter100|11364_ , \new_Sorter100|11365_ ,
    \new_Sorter100|11366_ , \new_Sorter100|11367_ , \new_Sorter100|11368_ ,
    \new_Sorter100|11369_ , \new_Sorter100|11370_ , \new_Sorter100|11371_ ,
    \new_Sorter100|11372_ , \new_Sorter100|11373_ , \new_Sorter100|11374_ ,
    \new_Sorter100|11375_ , \new_Sorter100|11376_ , \new_Sorter100|11377_ ,
    \new_Sorter100|11378_ , \new_Sorter100|11379_ , \new_Sorter100|11380_ ,
    \new_Sorter100|11381_ , \new_Sorter100|11382_ , \new_Sorter100|11383_ ,
    \new_Sorter100|11384_ , \new_Sorter100|11385_ , \new_Sorter100|11386_ ,
    \new_Sorter100|11387_ , \new_Sorter100|11388_ , \new_Sorter100|11389_ ,
    \new_Sorter100|11390_ , \new_Sorter100|11391_ , \new_Sorter100|11392_ ,
    \new_Sorter100|11393_ , \new_Sorter100|11394_ , \new_Sorter100|11395_ ,
    \new_Sorter100|11396_ , \new_Sorter100|11397_ , \new_Sorter100|11398_ ,
    \new_Sorter100|11400_ , \new_Sorter100|11401_ , \new_Sorter100|11402_ ,
    \new_Sorter100|11403_ , \new_Sorter100|11404_ , \new_Sorter100|11405_ ,
    \new_Sorter100|11406_ , \new_Sorter100|11407_ , \new_Sorter100|11408_ ,
    \new_Sorter100|11409_ , \new_Sorter100|11410_ , \new_Sorter100|11411_ ,
    \new_Sorter100|11412_ , \new_Sorter100|11413_ , \new_Sorter100|11414_ ,
    \new_Sorter100|11415_ , \new_Sorter100|11416_ , \new_Sorter100|11417_ ,
    \new_Sorter100|11418_ , \new_Sorter100|11419_ , \new_Sorter100|11420_ ,
    \new_Sorter100|11421_ , \new_Sorter100|11422_ , \new_Sorter100|11423_ ,
    \new_Sorter100|11424_ , \new_Sorter100|11425_ , \new_Sorter100|11426_ ,
    \new_Sorter100|11427_ , \new_Sorter100|11428_ , \new_Sorter100|11429_ ,
    \new_Sorter100|11430_ , \new_Sorter100|11431_ , \new_Sorter100|11432_ ,
    \new_Sorter100|11433_ , \new_Sorter100|11434_ , \new_Sorter100|11435_ ,
    \new_Sorter100|11436_ , \new_Sorter100|11437_ , \new_Sorter100|11438_ ,
    \new_Sorter100|11439_ , \new_Sorter100|11440_ , \new_Sorter100|11441_ ,
    \new_Sorter100|11442_ , \new_Sorter100|11443_ , \new_Sorter100|11444_ ,
    \new_Sorter100|11445_ , \new_Sorter100|11446_ , \new_Sorter100|11447_ ,
    \new_Sorter100|11448_ , \new_Sorter100|11449_ , \new_Sorter100|11450_ ,
    \new_Sorter100|11451_ , \new_Sorter100|11452_ , \new_Sorter100|11453_ ,
    \new_Sorter100|11454_ , \new_Sorter100|11455_ , \new_Sorter100|11456_ ,
    \new_Sorter100|11457_ , \new_Sorter100|11458_ , \new_Sorter100|11459_ ,
    \new_Sorter100|11460_ , \new_Sorter100|11461_ , \new_Sorter100|11462_ ,
    \new_Sorter100|11463_ , \new_Sorter100|11464_ , \new_Sorter100|11465_ ,
    \new_Sorter100|11466_ , \new_Sorter100|11467_ , \new_Sorter100|11468_ ,
    \new_Sorter100|11469_ , \new_Sorter100|11470_ , \new_Sorter100|11471_ ,
    \new_Sorter100|11472_ , \new_Sorter100|11473_ , \new_Sorter100|11474_ ,
    \new_Sorter100|11475_ , \new_Sorter100|11476_ , \new_Sorter100|11477_ ,
    \new_Sorter100|11478_ , \new_Sorter100|11479_ , \new_Sorter100|11480_ ,
    \new_Sorter100|11481_ , \new_Sorter100|11482_ , \new_Sorter100|11483_ ,
    \new_Sorter100|11484_ , \new_Sorter100|11485_ , \new_Sorter100|11486_ ,
    \new_Sorter100|11487_ , \new_Sorter100|11488_ , \new_Sorter100|11489_ ,
    \new_Sorter100|11490_ , \new_Sorter100|11491_ , \new_Sorter100|11492_ ,
    \new_Sorter100|11493_ , \new_Sorter100|11494_ , \new_Sorter100|11495_ ,
    \new_Sorter100|11496_ , \new_Sorter100|11497_ , \new_Sorter100|11498_ ,
    \new_Sorter100|11499_ , \new_Sorter100|11500_ , \new_Sorter100|11599_ ,
    \new_Sorter100|11501_ , \new_Sorter100|11502_ , \new_Sorter100|11503_ ,
    \new_Sorter100|11504_ , \new_Sorter100|11505_ , \new_Sorter100|11506_ ,
    \new_Sorter100|11507_ , \new_Sorter100|11508_ , \new_Sorter100|11509_ ,
    \new_Sorter100|11510_ , \new_Sorter100|11511_ , \new_Sorter100|11512_ ,
    \new_Sorter100|11513_ , \new_Sorter100|11514_ , \new_Sorter100|11515_ ,
    \new_Sorter100|11516_ , \new_Sorter100|11517_ , \new_Sorter100|11518_ ,
    \new_Sorter100|11519_ , \new_Sorter100|11520_ , \new_Sorter100|11521_ ,
    \new_Sorter100|11522_ , \new_Sorter100|11523_ , \new_Sorter100|11524_ ,
    \new_Sorter100|11525_ , \new_Sorter100|11526_ , \new_Sorter100|11527_ ,
    \new_Sorter100|11528_ , \new_Sorter100|11529_ , \new_Sorter100|11530_ ,
    \new_Sorter100|11531_ , \new_Sorter100|11532_ , \new_Sorter100|11533_ ,
    \new_Sorter100|11534_ , \new_Sorter100|11535_ , \new_Sorter100|11536_ ,
    \new_Sorter100|11537_ , \new_Sorter100|11538_ , \new_Sorter100|11539_ ,
    \new_Sorter100|11540_ , \new_Sorter100|11541_ , \new_Sorter100|11542_ ,
    \new_Sorter100|11543_ , \new_Sorter100|11544_ , \new_Sorter100|11545_ ,
    \new_Sorter100|11546_ , \new_Sorter100|11547_ , \new_Sorter100|11548_ ,
    \new_Sorter100|11549_ , \new_Sorter100|11550_ , \new_Sorter100|11551_ ,
    \new_Sorter100|11552_ , \new_Sorter100|11553_ , \new_Sorter100|11554_ ,
    \new_Sorter100|11555_ , \new_Sorter100|11556_ , \new_Sorter100|11557_ ,
    \new_Sorter100|11558_ , \new_Sorter100|11559_ , \new_Sorter100|11560_ ,
    \new_Sorter100|11561_ , \new_Sorter100|11562_ , \new_Sorter100|11563_ ,
    \new_Sorter100|11564_ , \new_Sorter100|11565_ , \new_Sorter100|11566_ ,
    \new_Sorter100|11567_ , \new_Sorter100|11568_ , \new_Sorter100|11569_ ,
    \new_Sorter100|11570_ , \new_Sorter100|11571_ , \new_Sorter100|11572_ ,
    \new_Sorter100|11573_ , \new_Sorter100|11574_ , \new_Sorter100|11575_ ,
    \new_Sorter100|11576_ , \new_Sorter100|11577_ , \new_Sorter100|11578_ ,
    \new_Sorter100|11579_ , \new_Sorter100|11580_ , \new_Sorter100|11581_ ,
    \new_Sorter100|11582_ , \new_Sorter100|11583_ , \new_Sorter100|11584_ ,
    \new_Sorter100|11585_ , \new_Sorter100|11586_ , \new_Sorter100|11587_ ,
    \new_Sorter100|11588_ , \new_Sorter100|11589_ , \new_Sorter100|11590_ ,
    \new_Sorter100|11591_ , \new_Sorter100|11592_ , \new_Sorter100|11593_ ,
    \new_Sorter100|11594_ , \new_Sorter100|11595_ , \new_Sorter100|11596_ ,
    \new_Sorter100|11597_ , \new_Sorter100|11598_ , \new_Sorter100|11600_ ,
    \new_Sorter100|11601_ , \new_Sorter100|11602_ , \new_Sorter100|11603_ ,
    \new_Sorter100|11604_ , \new_Sorter100|11605_ , \new_Sorter100|11606_ ,
    \new_Sorter100|11607_ , \new_Sorter100|11608_ , \new_Sorter100|11609_ ,
    \new_Sorter100|11610_ , \new_Sorter100|11611_ , \new_Sorter100|11612_ ,
    \new_Sorter100|11613_ , \new_Sorter100|11614_ , \new_Sorter100|11615_ ,
    \new_Sorter100|11616_ , \new_Sorter100|11617_ , \new_Sorter100|11618_ ,
    \new_Sorter100|11619_ , \new_Sorter100|11620_ , \new_Sorter100|11621_ ,
    \new_Sorter100|11622_ , \new_Sorter100|11623_ , \new_Sorter100|11624_ ,
    \new_Sorter100|11625_ , \new_Sorter100|11626_ , \new_Sorter100|11627_ ,
    \new_Sorter100|11628_ , \new_Sorter100|11629_ , \new_Sorter100|11630_ ,
    \new_Sorter100|11631_ , \new_Sorter100|11632_ , \new_Sorter100|11633_ ,
    \new_Sorter100|11634_ , \new_Sorter100|11635_ , \new_Sorter100|11636_ ,
    \new_Sorter100|11637_ , \new_Sorter100|11638_ , \new_Sorter100|11639_ ,
    \new_Sorter100|11640_ , \new_Sorter100|11641_ , \new_Sorter100|11642_ ,
    \new_Sorter100|11643_ , \new_Sorter100|11644_ , \new_Sorter100|11645_ ,
    \new_Sorter100|11646_ , \new_Sorter100|11647_ , \new_Sorter100|11648_ ,
    \new_Sorter100|11649_ , \new_Sorter100|11650_ , \new_Sorter100|11651_ ,
    \new_Sorter100|11652_ , \new_Sorter100|11653_ , \new_Sorter100|11654_ ,
    \new_Sorter100|11655_ , \new_Sorter100|11656_ , \new_Sorter100|11657_ ,
    \new_Sorter100|11658_ , \new_Sorter100|11659_ , \new_Sorter100|11660_ ,
    \new_Sorter100|11661_ , \new_Sorter100|11662_ , \new_Sorter100|11663_ ,
    \new_Sorter100|11664_ , \new_Sorter100|11665_ , \new_Sorter100|11666_ ,
    \new_Sorter100|11667_ , \new_Sorter100|11668_ , \new_Sorter100|11669_ ,
    \new_Sorter100|11670_ , \new_Sorter100|11671_ , \new_Sorter100|11672_ ,
    \new_Sorter100|11673_ , \new_Sorter100|11674_ , \new_Sorter100|11675_ ,
    \new_Sorter100|11676_ , \new_Sorter100|11677_ , \new_Sorter100|11678_ ,
    \new_Sorter100|11679_ , \new_Sorter100|11680_ , \new_Sorter100|11681_ ,
    \new_Sorter100|11682_ , \new_Sorter100|11683_ , \new_Sorter100|11684_ ,
    \new_Sorter100|11685_ , \new_Sorter100|11686_ , \new_Sorter100|11687_ ,
    \new_Sorter100|11688_ , \new_Sorter100|11689_ , \new_Sorter100|11690_ ,
    \new_Sorter100|11691_ , \new_Sorter100|11692_ , \new_Sorter100|11693_ ,
    \new_Sorter100|11694_ , \new_Sorter100|11695_ , \new_Sorter100|11696_ ,
    \new_Sorter100|11697_ , \new_Sorter100|11698_ , \new_Sorter100|11699_ ,
    \new_Sorter100|11700_ , \new_Sorter100|11799_ , \new_Sorter100|11701_ ,
    \new_Sorter100|11702_ , \new_Sorter100|11703_ , \new_Sorter100|11704_ ,
    \new_Sorter100|11705_ , \new_Sorter100|11706_ , \new_Sorter100|11707_ ,
    \new_Sorter100|11708_ , \new_Sorter100|11709_ , \new_Sorter100|11710_ ,
    \new_Sorter100|11711_ , \new_Sorter100|11712_ , \new_Sorter100|11713_ ,
    \new_Sorter100|11714_ , \new_Sorter100|11715_ , \new_Sorter100|11716_ ,
    \new_Sorter100|11717_ , \new_Sorter100|11718_ , \new_Sorter100|11719_ ,
    \new_Sorter100|11720_ , \new_Sorter100|11721_ , \new_Sorter100|11722_ ,
    \new_Sorter100|11723_ , \new_Sorter100|11724_ , \new_Sorter100|11725_ ,
    \new_Sorter100|11726_ , \new_Sorter100|11727_ , \new_Sorter100|11728_ ,
    \new_Sorter100|11729_ , \new_Sorter100|11730_ , \new_Sorter100|11731_ ,
    \new_Sorter100|11732_ , \new_Sorter100|11733_ , \new_Sorter100|11734_ ,
    \new_Sorter100|11735_ , \new_Sorter100|11736_ , \new_Sorter100|11737_ ,
    \new_Sorter100|11738_ , \new_Sorter100|11739_ , \new_Sorter100|11740_ ,
    \new_Sorter100|11741_ , \new_Sorter100|11742_ , \new_Sorter100|11743_ ,
    \new_Sorter100|11744_ , \new_Sorter100|11745_ , \new_Sorter100|11746_ ,
    \new_Sorter100|11747_ , \new_Sorter100|11748_ , \new_Sorter100|11749_ ,
    \new_Sorter100|11750_ , \new_Sorter100|11751_ , \new_Sorter100|11752_ ,
    \new_Sorter100|11753_ , \new_Sorter100|11754_ , \new_Sorter100|11755_ ,
    \new_Sorter100|11756_ , \new_Sorter100|11757_ , \new_Sorter100|11758_ ,
    \new_Sorter100|11759_ , \new_Sorter100|11760_ , \new_Sorter100|11761_ ,
    \new_Sorter100|11762_ , \new_Sorter100|11763_ , \new_Sorter100|11764_ ,
    \new_Sorter100|11765_ , \new_Sorter100|11766_ , \new_Sorter100|11767_ ,
    \new_Sorter100|11768_ , \new_Sorter100|11769_ , \new_Sorter100|11770_ ,
    \new_Sorter100|11771_ , \new_Sorter100|11772_ , \new_Sorter100|11773_ ,
    \new_Sorter100|11774_ , \new_Sorter100|11775_ , \new_Sorter100|11776_ ,
    \new_Sorter100|11777_ , \new_Sorter100|11778_ , \new_Sorter100|11779_ ,
    \new_Sorter100|11780_ , \new_Sorter100|11781_ , \new_Sorter100|11782_ ,
    \new_Sorter100|11783_ , \new_Sorter100|11784_ , \new_Sorter100|11785_ ,
    \new_Sorter100|11786_ , \new_Sorter100|11787_ , \new_Sorter100|11788_ ,
    \new_Sorter100|11789_ , \new_Sorter100|11790_ , \new_Sorter100|11791_ ,
    \new_Sorter100|11792_ , \new_Sorter100|11793_ , \new_Sorter100|11794_ ,
    \new_Sorter100|11795_ , \new_Sorter100|11796_ , \new_Sorter100|11797_ ,
    \new_Sorter100|11798_ , \new_Sorter100|11800_ , \new_Sorter100|11801_ ,
    \new_Sorter100|11802_ , \new_Sorter100|11803_ , \new_Sorter100|11804_ ,
    \new_Sorter100|11805_ , \new_Sorter100|11806_ , \new_Sorter100|11807_ ,
    \new_Sorter100|11808_ , \new_Sorter100|11809_ , \new_Sorter100|11810_ ,
    \new_Sorter100|11811_ , \new_Sorter100|11812_ , \new_Sorter100|11813_ ,
    \new_Sorter100|11814_ , \new_Sorter100|11815_ , \new_Sorter100|11816_ ,
    \new_Sorter100|11817_ , \new_Sorter100|11818_ , \new_Sorter100|11819_ ,
    \new_Sorter100|11820_ , \new_Sorter100|11821_ , \new_Sorter100|11822_ ,
    \new_Sorter100|11823_ , \new_Sorter100|11824_ , \new_Sorter100|11825_ ,
    \new_Sorter100|11826_ , \new_Sorter100|11827_ , \new_Sorter100|11828_ ,
    \new_Sorter100|11829_ , \new_Sorter100|11830_ , \new_Sorter100|11831_ ,
    \new_Sorter100|11832_ , \new_Sorter100|11833_ , \new_Sorter100|11834_ ,
    \new_Sorter100|11835_ , \new_Sorter100|11836_ , \new_Sorter100|11837_ ,
    \new_Sorter100|11838_ , \new_Sorter100|11839_ , \new_Sorter100|11840_ ,
    \new_Sorter100|11841_ , \new_Sorter100|11842_ , \new_Sorter100|11843_ ,
    \new_Sorter100|11844_ , \new_Sorter100|11845_ , \new_Sorter100|11846_ ,
    \new_Sorter100|11847_ , \new_Sorter100|11848_ , \new_Sorter100|11849_ ,
    \new_Sorter100|11850_ , \new_Sorter100|11851_ , \new_Sorter100|11852_ ,
    \new_Sorter100|11853_ , \new_Sorter100|11854_ , \new_Sorter100|11855_ ,
    \new_Sorter100|11856_ , \new_Sorter100|11857_ , \new_Sorter100|11858_ ,
    \new_Sorter100|11859_ , \new_Sorter100|11860_ , \new_Sorter100|11861_ ,
    \new_Sorter100|11862_ , \new_Sorter100|11863_ , \new_Sorter100|11864_ ,
    \new_Sorter100|11865_ , \new_Sorter100|11866_ , \new_Sorter100|11867_ ,
    \new_Sorter100|11868_ , \new_Sorter100|11869_ , \new_Sorter100|11870_ ,
    \new_Sorter100|11871_ , \new_Sorter100|11872_ , \new_Sorter100|11873_ ,
    \new_Sorter100|11874_ , \new_Sorter100|11875_ , \new_Sorter100|11876_ ,
    \new_Sorter100|11877_ , \new_Sorter100|11878_ , \new_Sorter100|11879_ ,
    \new_Sorter100|11880_ , \new_Sorter100|11881_ , \new_Sorter100|11882_ ,
    \new_Sorter100|11883_ , \new_Sorter100|11884_ , \new_Sorter100|11885_ ,
    \new_Sorter100|11886_ , \new_Sorter100|11887_ , \new_Sorter100|11888_ ,
    \new_Sorter100|11889_ , \new_Sorter100|11890_ , \new_Sorter100|11891_ ,
    \new_Sorter100|11892_ , \new_Sorter100|11893_ , \new_Sorter100|11894_ ,
    \new_Sorter100|11895_ , \new_Sorter100|11896_ , \new_Sorter100|11897_ ,
    \new_Sorter100|11898_ , \new_Sorter100|11899_ , \new_Sorter100|11900_ ,
    \new_Sorter100|11999_ , \new_Sorter100|11901_ , \new_Sorter100|11902_ ,
    \new_Sorter100|11903_ , \new_Sorter100|11904_ , \new_Sorter100|11905_ ,
    \new_Sorter100|11906_ , \new_Sorter100|11907_ , \new_Sorter100|11908_ ,
    \new_Sorter100|11909_ , \new_Sorter100|11910_ , \new_Sorter100|11911_ ,
    \new_Sorter100|11912_ , \new_Sorter100|11913_ , \new_Sorter100|11914_ ,
    \new_Sorter100|11915_ , \new_Sorter100|11916_ , \new_Sorter100|11917_ ,
    \new_Sorter100|11918_ , \new_Sorter100|11919_ , \new_Sorter100|11920_ ,
    \new_Sorter100|11921_ , \new_Sorter100|11922_ , \new_Sorter100|11923_ ,
    \new_Sorter100|11924_ , \new_Sorter100|11925_ , \new_Sorter100|11926_ ,
    \new_Sorter100|11927_ , \new_Sorter100|11928_ , \new_Sorter100|11929_ ,
    \new_Sorter100|11930_ , \new_Sorter100|11931_ , \new_Sorter100|11932_ ,
    \new_Sorter100|11933_ , \new_Sorter100|11934_ , \new_Sorter100|11935_ ,
    \new_Sorter100|11936_ , \new_Sorter100|11937_ , \new_Sorter100|11938_ ,
    \new_Sorter100|11939_ , \new_Sorter100|11940_ , \new_Sorter100|11941_ ,
    \new_Sorter100|11942_ , \new_Sorter100|11943_ , \new_Sorter100|11944_ ,
    \new_Sorter100|11945_ , \new_Sorter100|11946_ , \new_Sorter100|11947_ ,
    \new_Sorter100|11948_ , \new_Sorter100|11949_ , \new_Sorter100|11950_ ,
    \new_Sorter100|11951_ , \new_Sorter100|11952_ , \new_Sorter100|11953_ ,
    \new_Sorter100|11954_ , \new_Sorter100|11955_ , \new_Sorter100|11956_ ,
    \new_Sorter100|11957_ , \new_Sorter100|11958_ , \new_Sorter100|11959_ ,
    \new_Sorter100|11960_ , \new_Sorter100|11961_ , \new_Sorter100|11962_ ,
    \new_Sorter100|11963_ , \new_Sorter100|11964_ , \new_Sorter100|11965_ ,
    \new_Sorter100|11966_ , \new_Sorter100|11967_ , \new_Sorter100|11968_ ,
    \new_Sorter100|11969_ , \new_Sorter100|11970_ , \new_Sorter100|11971_ ,
    \new_Sorter100|11972_ , \new_Sorter100|11973_ , \new_Sorter100|11974_ ,
    \new_Sorter100|11975_ , \new_Sorter100|11976_ , \new_Sorter100|11977_ ,
    \new_Sorter100|11978_ , \new_Sorter100|11979_ , \new_Sorter100|11980_ ,
    \new_Sorter100|11981_ , \new_Sorter100|11982_ , \new_Sorter100|11983_ ,
    \new_Sorter100|11984_ , \new_Sorter100|11985_ , \new_Sorter100|11986_ ,
    \new_Sorter100|11987_ , \new_Sorter100|11988_ , \new_Sorter100|11989_ ,
    \new_Sorter100|11990_ , \new_Sorter100|11991_ , \new_Sorter100|11992_ ,
    \new_Sorter100|11993_ , \new_Sorter100|11994_ , \new_Sorter100|11995_ ,
    \new_Sorter100|11996_ , \new_Sorter100|11997_ , \new_Sorter100|11998_ ,
    \new_Sorter100|12000_ , \new_Sorter100|12001_ , \new_Sorter100|12002_ ,
    \new_Sorter100|12003_ , \new_Sorter100|12004_ , \new_Sorter100|12005_ ,
    \new_Sorter100|12006_ , \new_Sorter100|12007_ , \new_Sorter100|12008_ ,
    \new_Sorter100|12009_ , \new_Sorter100|12010_ , \new_Sorter100|12011_ ,
    \new_Sorter100|12012_ , \new_Sorter100|12013_ , \new_Sorter100|12014_ ,
    \new_Sorter100|12015_ , \new_Sorter100|12016_ , \new_Sorter100|12017_ ,
    \new_Sorter100|12018_ , \new_Sorter100|12019_ , \new_Sorter100|12020_ ,
    \new_Sorter100|12021_ , \new_Sorter100|12022_ , \new_Sorter100|12023_ ,
    \new_Sorter100|12024_ , \new_Sorter100|12025_ , \new_Sorter100|12026_ ,
    \new_Sorter100|12027_ , \new_Sorter100|12028_ , \new_Sorter100|12029_ ,
    \new_Sorter100|12030_ , \new_Sorter100|12031_ , \new_Sorter100|12032_ ,
    \new_Sorter100|12033_ , \new_Sorter100|12034_ , \new_Sorter100|12035_ ,
    \new_Sorter100|12036_ , \new_Sorter100|12037_ , \new_Sorter100|12038_ ,
    \new_Sorter100|12039_ , \new_Sorter100|12040_ , \new_Sorter100|12041_ ,
    \new_Sorter100|12042_ , \new_Sorter100|12043_ , \new_Sorter100|12044_ ,
    \new_Sorter100|12045_ , \new_Sorter100|12046_ , \new_Sorter100|12047_ ,
    \new_Sorter100|12048_ , \new_Sorter100|12049_ , \new_Sorter100|12050_ ,
    \new_Sorter100|12051_ , \new_Sorter100|12052_ , \new_Sorter100|12053_ ,
    \new_Sorter100|12054_ , \new_Sorter100|12055_ , \new_Sorter100|12056_ ,
    \new_Sorter100|12057_ , \new_Sorter100|12058_ , \new_Sorter100|12059_ ,
    \new_Sorter100|12060_ , \new_Sorter100|12061_ , \new_Sorter100|12062_ ,
    \new_Sorter100|12063_ , \new_Sorter100|12064_ , \new_Sorter100|12065_ ,
    \new_Sorter100|12066_ , \new_Sorter100|12067_ , \new_Sorter100|12068_ ,
    \new_Sorter100|12069_ , \new_Sorter100|12070_ , \new_Sorter100|12071_ ,
    \new_Sorter100|12072_ , \new_Sorter100|12073_ , \new_Sorter100|12074_ ,
    \new_Sorter100|12075_ , \new_Sorter100|12076_ , \new_Sorter100|12077_ ,
    \new_Sorter100|12078_ , \new_Sorter100|12079_ , \new_Sorter100|12080_ ,
    \new_Sorter100|12081_ , \new_Sorter100|12082_ , \new_Sorter100|12083_ ,
    \new_Sorter100|12084_ , \new_Sorter100|12085_ , \new_Sorter100|12086_ ,
    \new_Sorter100|12087_ , \new_Sorter100|12088_ , \new_Sorter100|12089_ ,
    \new_Sorter100|12090_ , \new_Sorter100|12091_ , \new_Sorter100|12092_ ,
    \new_Sorter100|12093_ , \new_Sorter100|12094_ , \new_Sorter100|12095_ ,
    \new_Sorter100|12096_ , \new_Sorter100|12097_ , \new_Sorter100|12098_ ,
    \new_Sorter100|12099_ , \new_Sorter100|12100_ , \new_Sorter100|12199_ ,
    \new_Sorter100|12101_ , \new_Sorter100|12102_ , \new_Sorter100|12103_ ,
    \new_Sorter100|12104_ , \new_Sorter100|12105_ , \new_Sorter100|12106_ ,
    \new_Sorter100|12107_ , \new_Sorter100|12108_ , \new_Sorter100|12109_ ,
    \new_Sorter100|12110_ , \new_Sorter100|12111_ , \new_Sorter100|12112_ ,
    \new_Sorter100|12113_ , \new_Sorter100|12114_ , \new_Sorter100|12115_ ,
    \new_Sorter100|12116_ , \new_Sorter100|12117_ , \new_Sorter100|12118_ ,
    \new_Sorter100|12119_ , \new_Sorter100|12120_ , \new_Sorter100|12121_ ,
    \new_Sorter100|12122_ , \new_Sorter100|12123_ , \new_Sorter100|12124_ ,
    \new_Sorter100|12125_ , \new_Sorter100|12126_ , \new_Sorter100|12127_ ,
    \new_Sorter100|12128_ , \new_Sorter100|12129_ , \new_Sorter100|12130_ ,
    \new_Sorter100|12131_ , \new_Sorter100|12132_ , \new_Sorter100|12133_ ,
    \new_Sorter100|12134_ , \new_Sorter100|12135_ , \new_Sorter100|12136_ ,
    \new_Sorter100|12137_ , \new_Sorter100|12138_ , \new_Sorter100|12139_ ,
    \new_Sorter100|12140_ , \new_Sorter100|12141_ , \new_Sorter100|12142_ ,
    \new_Sorter100|12143_ , \new_Sorter100|12144_ , \new_Sorter100|12145_ ,
    \new_Sorter100|12146_ , \new_Sorter100|12147_ , \new_Sorter100|12148_ ,
    \new_Sorter100|12149_ , \new_Sorter100|12150_ , \new_Sorter100|12151_ ,
    \new_Sorter100|12152_ , \new_Sorter100|12153_ , \new_Sorter100|12154_ ,
    \new_Sorter100|12155_ , \new_Sorter100|12156_ , \new_Sorter100|12157_ ,
    \new_Sorter100|12158_ , \new_Sorter100|12159_ , \new_Sorter100|12160_ ,
    \new_Sorter100|12161_ , \new_Sorter100|12162_ , \new_Sorter100|12163_ ,
    \new_Sorter100|12164_ , \new_Sorter100|12165_ , \new_Sorter100|12166_ ,
    \new_Sorter100|12167_ , \new_Sorter100|12168_ , \new_Sorter100|12169_ ,
    \new_Sorter100|12170_ , \new_Sorter100|12171_ , \new_Sorter100|12172_ ,
    \new_Sorter100|12173_ , \new_Sorter100|12174_ , \new_Sorter100|12175_ ,
    \new_Sorter100|12176_ , \new_Sorter100|12177_ , \new_Sorter100|12178_ ,
    \new_Sorter100|12179_ , \new_Sorter100|12180_ , \new_Sorter100|12181_ ,
    \new_Sorter100|12182_ , \new_Sorter100|12183_ , \new_Sorter100|12184_ ,
    \new_Sorter100|12185_ , \new_Sorter100|12186_ , \new_Sorter100|12187_ ,
    \new_Sorter100|12188_ , \new_Sorter100|12189_ , \new_Sorter100|12190_ ,
    \new_Sorter100|12191_ , \new_Sorter100|12192_ , \new_Sorter100|12193_ ,
    \new_Sorter100|12194_ , \new_Sorter100|12195_ , \new_Sorter100|12196_ ,
    \new_Sorter100|12197_ , \new_Sorter100|12198_ , \new_Sorter100|12200_ ,
    \new_Sorter100|12201_ , \new_Sorter100|12202_ , \new_Sorter100|12203_ ,
    \new_Sorter100|12204_ , \new_Sorter100|12205_ , \new_Sorter100|12206_ ,
    \new_Sorter100|12207_ , \new_Sorter100|12208_ , \new_Sorter100|12209_ ,
    \new_Sorter100|12210_ , \new_Sorter100|12211_ , \new_Sorter100|12212_ ,
    \new_Sorter100|12213_ , \new_Sorter100|12214_ , \new_Sorter100|12215_ ,
    \new_Sorter100|12216_ , \new_Sorter100|12217_ , \new_Sorter100|12218_ ,
    \new_Sorter100|12219_ , \new_Sorter100|12220_ , \new_Sorter100|12221_ ,
    \new_Sorter100|12222_ , \new_Sorter100|12223_ , \new_Sorter100|12224_ ,
    \new_Sorter100|12225_ , \new_Sorter100|12226_ , \new_Sorter100|12227_ ,
    \new_Sorter100|12228_ , \new_Sorter100|12229_ , \new_Sorter100|12230_ ,
    \new_Sorter100|12231_ , \new_Sorter100|12232_ , \new_Sorter100|12233_ ,
    \new_Sorter100|12234_ , \new_Sorter100|12235_ , \new_Sorter100|12236_ ,
    \new_Sorter100|12237_ , \new_Sorter100|12238_ , \new_Sorter100|12239_ ,
    \new_Sorter100|12240_ , \new_Sorter100|12241_ , \new_Sorter100|12242_ ,
    \new_Sorter100|12243_ , \new_Sorter100|12244_ , \new_Sorter100|12245_ ,
    \new_Sorter100|12246_ , \new_Sorter100|12247_ , \new_Sorter100|12248_ ,
    \new_Sorter100|12249_ , \new_Sorter100|12250_ , \new_Sorter100|12251_ ,
    \new_Sorter100|12252_ , \new_Sorter100|12253_ , \new_Sorter100|12254_ ,
    \new_Sorter100|12255_ , \new_Sorter100|12256_ , \new_Sorter100|12257_ ,
    \new_Sorter100|12258_ , \new_Sorter100|12259_ , \new_Sorter100|12260_ ,
    \new_Sorter100|12261_ , \new_Sorter100|12262_ , \new_Sorter100|12263_ ,
    \new_Sorter100|12264_ , \new_Sorter100|12265_ , \new_Sorter100|12266_ ,
    \new_Sorter100|12267_ , \new_Sorter100|12268_ , \new_Sorter100|12269_ ,
    \new_Sorter100|12270_ , \new_Sorter100|12271_ , \new_Sorter100|12272_ ,
    \new_Sorter100|12273_ , \new_Sorter100|12274_ , \new_Sorter100|12275_ ,
    \new_Sorter100|12276_ , \new_Sorter100|12277_ , \new_Sorter100|12278_ ,
    \new_Sorter100|12279_ , \new_Sorter100|12280_ , \new_Sorter100|12281_ ,
    \new_Sorter100|12282_ , \new_Sorter100|12283_ , \new_Sorter100|12284_ ,
    \new_Sorter100|12285_ , \new_Sorter100|12286_ , \new_Sorter100|12287_ ,
    \new_Sorter100|12288_ , \new_Sorter100|12289_ , \new_Sorter100|12290_ ,
    \new_Sorter100|12291_ , \new_Sorter100|12292_ , \new_Sorter100|12293_ ,
    \new_Sorter100|12294_ , \new_Sorter100|12295_ , \new_Sorter100|12296_ ,
    \new_Sorter100|12297_ , \new_Sorter100|12298_ , \new_Sorter100|12299_ ,
    \new_Sorter100|12300_ , \new_Sorter100|12399_ , \new_Sorter100|12301_ ,
    \new_Sorter100|12302_ , \new_Sorter100|12303_ , \new_Sorter100|12304_ ,
    \new_Sorter100|12305_ , \new_Sorter100|12306_ , \new_Sorter100|12307_ ,
    \new_Sorter100|12308_ , \new_Sorter100|12309_ , \new_Sorter100|12310_ ,
    \new_Sorter100|12311_ , \new_Sorter100|12312_ , \new_Sorter100|12313_ ,
    \new_Sorter100|12314_ , \new_Sorter100|12315_ , \new_Sorter100|12316_ ,
    \new_Sorter100|12317_ , \new_Sorter100|12318_ , \new_Sorter100|12319_ ,
    \new_Sorter100|12320_ , \new_Sorter100|12321_ , \new_Sorter100|12322_ ,
    \new_Sorter100|12323_ , \new_Sorter100|12324_ , \new_Sorter100|12325_ ,
    \new_Sorter100|12326_ , \new_Sorter100|12327_ , \new_Sorter100|12328_ ,
    \new_Sorter100|12329_ , \new_Sorter100|12330_ , \new_Sorter100|12331_ ,
    \new_Sorter100|12332_ , \new_Sorter100|12333_ , \new_Sorter100|12334_ ,
    \new_Sorter100|12335_ , \new_Sorter100|12336_ , \new_Sorter100|12337_ ,
    \new_Sorter100|12338_ , \new_Sorter100|12339_ , \new_Sorter100|12340_ ,
    \new_Sorter100|12341_ , \new_Sorter100|12342_ , \new_Sorter100|12343_ ,
    \new_Sorter100|12344_ , \new_Sorter100|12345_ , \new_Sorter100|12346_ ,
    \new_Sorter100|12347_ , \new_Sorter100|12348_ , \new_Sorter100|12349_ ,
    \new_Sorter100|12350_ , \new_Sorter100|12351_ , \new_Sorter100|12352_ ,
    \new_Sorter100|12353_ , \new_Sorter100|12354_ , \new_Sorter100|12355_ ,
    \new_Sorter100|12356_ , \new_Sorter100|12357_ , \new_Sorter100|12358_ ,
    \new_Sorter100|12359_ , \new_Sorter100|12360_ , \new_Sorter100|12361_ ,
    \new_Sorter100|12362_ , \new_Sorter100|12363_ , \new_Sorter100|12364_ ,
    \new_Sorter100|12365_ , \new_Sorter100|12366_ , \new_Sorter100|12367_ ,
    \new_Sorter100|12368_ , \new_Sorter100|12369_ , \new_Sorter100|12370_ ,
    \new_Sorter100|12371_ , \new_Sorter100|12372_ , \new_Sorter100|12373_ ,
    \new_Sorter100|12374_ , \new_Sorter100|12375_ , \new_Sorter100|12376_ ,
    \new_Sorter100|12377_ , \new_Sorter100|12378_ , \new_Sorter100|12379_ ,
    \new_Sorter100|12380_ , \new_Sorter100|12381_ , \new_Sorter100|12382_ ,
    \new_Sorter100|12383_ , \new_Sorter100|12384_ , \new_Sorter100|12385_ ,
    \new_Sorter100|12386_ , \new_Sorter100|12387_ , \new_Sorter100|12388_ ,
    \new_Sorter100|12389_ , \new_Sorter100|12390_ , \new_Sorter100|12391_ ,
    \new_Sorter100|12392_ , \new_Sorter100|12393_ , \new_Sorter100|12394_ ,
    \new_Sorter100|12395_ , \new_Sorter100|12396_ , \new_Sorter100|12397_ ,
    \new_Sorter100|12398_ , \new_Sorter100|12400_ , \new_Sorter100|12401_ ,
    \new_Sorter100|12402_ , \new_Sorter100|12403_ , \new_Sorter100|12404_ ,
    \new_Sorter100|12405_ , \new_Sorter100|12406_ , \new_Sorter100|12407_ ,
    \new_Sorter100|12408_ , \new_Sorter100|12409_ , \new_Sorter100|12410_ ,
    \new_Sorter100|12411_ , \new_Sorter100|12412_ , \new_Sorter100|12413_ ,
    \new_Sorter100|12414_ , \new_Sorter100|12415_ , \new_Sorter100|12416_ ,
    \new_Sorter100|12417_ , \new_Sorter100|12418_ , \new_Sorter100|12419_ ,
    \new_Sorter100|12420_ , \new_Sorter100|12421_ , \new_Sorter100|12422_ ,
    \new_Sorter100|12423_ , \new_Sorter100|12424_ , \new_Sorter100|12425_ ,
    \new_Sorter100|12426_ , \new_Sorter100|12427_ , \new_Sorter100|12428_ ,
    \new_Sorter100|12429_ , \new_Sorter100|12430_ , \new_Sorter100|12431_ ,
    \new_Sorter100|12432_ , \new_Sorter100|12433_ , \new_Sorter100|12434_ ,
    \new_Sorter100|12435_ , \new_Sorter100|12436_ , \new_Sorter100|12437_ ,
    \new_Sorter100|12438_ , \new_Sorter100|12439_ , \new_Sorter100|12440_ ,
    \new_Sorter100|12441_ , \new_Sorter100|12442_ , \new_Sorter100|12443_ ,
    \new_Sorter100|12444_ , \new_Sorter100|12445_ , \new_Sorter100|12446_ ,
    \new_Sorter100|12447_ , \new_Sorter100|12448_ , \new_Sorter100|12449_ ,
    \new_Sorter100|12450_ , \new_Sorter100|12451_ , \new_Sorter100|12452_ ,
    \new_Sorter100|12453_ , \new_Sorter100|12454_ , \new_Sorter100|12455_ ,
    \new_Sorter100|12456_ , \new_Sorter100|12457_ , \new_Sorter100|12458_ ,
    \new_Sorter100|12459_ , \new_Sorter100|12460_ , \new_Sorter100|12461_ ,
    \new_Sorter100|12462_ , \new_Sorter100|12463_ , \new_Sorter100|12464_ ,
    \new_Sorter100|12465_ , \new_Sorter100|12466_ , \new_Sorter100|12467_ ,
    \new_Sorter100|12468_ , \new_Sorter100|12469_ , \new_Sorter100|12470_ ,
    \new_Sorter100|12471_ , \new_Sorter100|12472_ , \new_Sorter100|12473_ ,
    \new_Sorter100|12474_ , \new_Sorter100|12475_ , \new_Sorter100|12476_ ,
    \new_Sorter100|12477_ , \new_Sorter100|12478_ , \new_Sorter100|12479_ ,
    \new_Sorter100|12480_ , \new_Sorter100|12481_ , \new_Sorter100|12482_ ,
    \new_Sorter100|12483_ , \new_Sorter100|12484_ , \new_Sorter100|12485_ ,
    \new_Sorter100|12486_ , \new_Sorter100|12487_ , \new_Sorter100|12488_ ,
    \new_Sorter100|12489_ , \new_Sorter100|12490_ , \new_Sorter100|12491_ ,
    \new_Sorter100|12492_ , \new_Sorter100|12493_ , \new_Sorter100|12494_ ,
    \new_Sorter100|12495_ , \new_Sorter100|12496_ , \new_Sorter100|12497_ ,
    \new_Sorter100|12498_ , \new_Sorter100|12499_ , \new_Sorter100|12500_ ,
    \new_Sorter100|12599_ , \new_Sorter100|12501_ , \new_Sorter100|12502_ ,
    \new_Sorter100|12503_ , \new_Sorter100|12504_ , \new_Sorter100|12505_ ,
    \new_Sorter100|12506_ , \new_Sorter100|12507_ , \new_Sorter100|12508_ ,
    \new_Sorter100|12509_ , \new_Sorter100|12510_ , \new_Sorter100|12511_ ,
    \new_Sorter100|12512_ , \new_Sorter100|12513_ , \new_Sorter100|12514_ ,
    \new_Sorter100|12515_ , \new_Sorter100|12516_ , \new_Sorter100|12517_ ,
    \new_Sorter100|12518_ , \new_Sorter100|12519_ , \new_Sorter100|12520_ ,
    \new_Sorter100|12521_ , \new_Sorter100|12522_ , \new_Sorter100|12523_ ,
    \new_Sorter100|12524_ , \new_Sorter100|12525_ , \new_Sorter100|12526_ ,
    \new_Sorter100|12527_ , \new_Sorter100|12528_ , \new_Sorter100|12529_ ,
    \new_Sorter100|12530_ , \new_Sorter100|12531_ , \new_Sorter100|12532_ ,
    \new_Sorter100|12533_ , \new_Sorter100|12534_ , \new_Sorter100|12535_ ,
    \new_Sorter100|12536_ , \new_Sorter100|12537_ , \new_Sorter100|12538_ ,
    \new_Sorter100|12539_ , \new_Sorter100|12540_ , \new_Sorter100|12541_ ,
    \new_Sorter100|12542_ , \new_Sorter100|12543_ , \new_Sorter100|12544_ ,
    \new_Sorter100|12545_ , \new_Sorter100|12546_ , \new_Sorter100|12547_ ,
    \new_Sorter100|12548_ , \new_Sorter100|12549_ , \new_Sorter100|12550_ ,
    \new_Sorter100|12551_ , \new_Sorter100|12552_ , \new_Sorter100|12553_ ,
    \new_Sorter100|12554_ , \new_Sorter100|12555_ , \new_Sorter100|12556_ ,
    \new_Sorter100|12557_ , \new_Sorter100|12558_ , \new_Sorter100|12559_ ,
    \new_Sorter100|12560_ , \new_Sorter100|12561_ , \new_Sorter100|12562_ ,
    \new_Sorter100|12563_ , \new_Sorter100|12564_ , \new_Sorter100|12565_ ,
    \new_Sorter100|12566_ , \new_Sorter100|12567_ , \new_Sorter100|12568_ ,
    \new_Sorter100|12569_ , \new_Sorter100|12570_ , \new_Sorter100|12571_ ,
    \new_Sorter100|12572_ , \new_Sorter100|12573_ , \new_Sorter100|12574_ ,
    \new_Sorter100|12575_ , \new_Sorter100|12576_ , \new_Sorter100|12577_ ,
    \new_Sorter100|12578_ , \new_Sorter100|12579_ , \new_Sorter100|12580_ ,
    \new_Sorter100|12581_ , \new_Sorter100|12582_ , \new_Sorter100|12583_ ,
    \new_Sorter100|12584_ , \new_Sorter100|12585_ , \new_Sorter100|12586_ ,
    \new_Sorter100|12587_ , \new_Sorter100|12588_ , \new_Sorter100|12589_ ,
    \new_Sorter100|12590_ , \new_Sorter100|12591_ , \new_Sorter100|12592_ ,
    \new_Sorter100|12593_ , \new_Sorter100|12594_ , \new_Sorter100|12595_ ,
    \new_Sorter100|12596_ , \new_Sorter100|12597_ , \new_Sorter100|12598_ ,
    \new_Sorter100|12600_ , \new_Sorter100|12601_ , \new_Sorter100|12602_ ,
    \new_Sorter100|12603_ , \new_Sorter100|12604_ , \new_Sorter100|12605_ ,
    \new_Sorter100|12606_ , \new_Sorter100|12607_ , \new_Sorter100|12608_ ,
    \new_Sorter100|12609_ , \new_Sorter100|12610_ , \new_Sorter100|12611_ ,
    \new_Sorter100|12612_ , \new_Sorter100|12613_ , \new_Sorter100|12614_ ,
    \new_Sorter100|12615_ , \new_Sorter100|12616_ , \new_Sorter100|12617_ ,
    \new_Sorter100|12618_ , \new_Sorter100|12619_ , \new_Sorter100|12620_ ,
    \new_Sorter100|12621_ , \new_Sorter100|12622_ , \new_Sorter100|12623_ ,
    \new_Sorter100|12624_ , \new_Sorter100|12625_ , \new_Sorter100|12626_ ,
    \new_Sorter100|12627_ , \new_Sorter100|12628_ , \new_Sorter100|12629_ ,
    \new_Sorter100|12630_ , \new_Sorter100|12631_ , \new_Sorter100|12632_ ,
    \new_Sorter100|12633_ , \new_Sorter100|12634_ , \new_Sorter100|12635_ ,
    \new_Sorter100|12636_ , \new_Sorter100|12637_ , \new_Sorter100|12638_ ,
    \new_Sorter100|12639_ , \new_Sorter100|12640_ , \new_Sorter100|12641_ ,
    \new_Sorter100|12642_ , \new_Sorter100|12643_ , \new_Sorter100|12644_ ,
    \new_Sorter100|12645_ , \new_Sorter100|12646_ , \new_Sorter100|12647_ ,
    \new_Sorter100|12648_ , \new_Sorter100|12649_ , \new_Sorter100|12650_ ,
    \new_Sorter100|12651_ , \new_Sorter100|12652_ , \new_Sorter100|12653_ ,
    \new_Sorter100|12654_ , \new_Sorter100|12655_ , \new_Sorter100|12656_ ,
    \new_Sorter100|12657_ , \new_Sorter100|12658_ , \new_Sorter100|12659_ ,
    \new_Sorter100|12660_ , \new_Sorter100|12661_ , \new_Sorter100|12662_ ,
    \new_Sorter100|12663_ , \new_Sorter100|12664_ , \new_Sorter100|12665_ ,
    \new_Sorter100|12666_ , \new_Sorter100|12667_ , \new_Sorter100|12668_ ,
    \new_Sorter100|12669_ , \new_Sorter100|12670_ , \new_Sorter100|12671_ ,
    \new_Sorter100|12672_ , \new_Sorter100|12673_ , \new_Sorter100|12674_ ,
    \new_Sorter100|12675_ , \new_Sorter100|12676_ , \new_Sorter100|12677_ ,
    \new_Sorter100|12678_ , \new_Sorter100|12679_ , \new_Sorter100|12680_ ,
    \new_Sorter100|12681_ , \new_Sorter100|12682_ , \new_Sorter100|12683_ ,
    \new_Sorter100|12684_ , \new_Sorter100|12685_ , \new_Sorter100|12686_ ,
    \new_Sorter100|12687_ , \new_Sorter100|12688_ , \new_Sorter100|12689_ ,
    \new_Sorter100|12690_ , \new_Sorter100|12691_ , \new_Sorter100|12692_ ,
    \new_Sorter100|12693_ , \new_Sorter100|12694_ , \new_Sorter100|12695_ ,
    \new_Sorter100|12696_ , \new_Sorter100|12697_ , \new_Sorter100|12698_ ,
    \new_Sorter100|12699_ , \new_Sorter100|12700_ , \new_Sorter100|12799_ ,
    \new_Sorter100|12701_ , \new_Sorter100|12702_ , \new_Sorter100|12703_ ,
    \new_Sorter100|12704_ , \new_Sorter100|12705_ , \new_Sorter100|12706_ ,
    \new_Sorter100|12707_ , \new_Sorter100|12708_ , \new_Sorter100|12709_ ,
    \new_Sorter100|12710_ , \new_Sorter100|12711_ , \new_Sorter100|12712_ ,
    \new_Sorter100|12713_ , \new_Sorter100|12714_ , \new_Sorter100|12715_ ,
    \new_Sorter100|12716_ , \new_Sorter100|12717_ , \new_Sorter100|12718_ ,
    \new_Sorter100|12719_ , \new_Sorter100|12720_ , \new_Sorter100|12721_ ,
    \new_Sorter100|12722_ , \new_Sorter100|12723_ , \new_Sorter100|12724_ ,
    \new_Sorter100|12725_ , \new_Sorter100|12726_ , \new_Sorter100|12727_ ,
    \new_Sorter100|12728_ , \new_Sorter100|12729_ , \new_Sorter100|12730_ ,
    \new_Sorter100|12731_ , \new_Sorter100|12732_ , \new_Sorter100|12733_ ,
    \new_Sorter100|12734_ , \new_Sorter100|12735_ , \new_Sorter100|12736_ ,
    \new_Sorter100|12737_ , \new_Sorter100|12738_ , \new_Sorter100|12739_ ,
    \new_Sorter100|12740_ , \new_Sorter100|12741_ , \new_Sorter100|12742_ ,
    \new_Sorter100|12743_ , \new_Sorter100|12744_ , \new_Sorter100|12745_ ,
    \new_Sorter100|12746_ , \new_Sorter100|12747_ , \new_Sorter100|12748_ ,
    \new_Sorter100|12749_ , \new_Sorter100|12750_ , \new_Sorter100|12751_ ,
    \new_Sorter100|12752_ , \new_Sorter100|12753_ , \new_Sorter100|12754_ ,
    \new_Sorter100|12755_ , \new_Sorter100|12756_ , \new_Sorter100|12757_ ,
    \new_Sorter100|12758_ , \new_Sorter100|12759_ , \new_Sorter100|12760_ ,
    \new_Sorter100|12761_ , \new_Sorter100|12762_ , \new_Sorter100|12763_ ,
    \new_Sorter100|12764_ , \new_Sorter100|12765_ , \new_Sorter100|12766_ ,
    \new_Sorter100|12767_ , \new_Sorter100|12768_ , \new_Sorter100|12769_ ,
    \new_Sorter100|12770_ , \new_Sorter100|12771_ , \new_Sorter100|12772_ ,
    \new_Sorter100|12773_ , \new_Sorter100|12774_ , \new_Sorter100|12775_ ,
    \new_Sorter100|12776_ , \new_Sorter100|12777_ , \new_Sorter100|12778_ ,
    \new_Sorter100|12779_ , \new_Sorter100|12780_ , \new_Sorter100|12781_ ,
    \new_Sorter100|12782_ , \new_Sorter100|12783_ , \new_Sorter100|12784_ ,
    \new_Sorter100|12785_ , \new_Sorter100|12786_ , \new_Sorter100|12787_ ,
    \new_Sorter100|12788_ , \new_Sorter100|12789_ , \new_Sorter100|12790_ ,
    \new_Sorter100|12791_ , \new_Sorter100|12792_ , \new_Sorter100|12793_ ,
    \new_Sorter100|12794_ , \new_Sorter100|12795_ , \new_Sorter100|12796_ ,
    \new_Sorter100|12797_ , \new_Sorter100|12798_ , \new_Sorter100|12800_ ,
    \new_Sorter100|12801_ , \new_Sorter100|12802_ , \new_Sorter100|12803_ ,
    \new_Sorter100|12804_ , \new_Sorter100|12805_ , \new_Sorter100|12806_ ,
    \new_Sorter100|12807_ , \new_Sorter100|12808_ , \new_Sorter100|12809_ ,
    \new_Sorter100|12810_ , \new_Sorter100|12811_ , \new_Sorter100|12812_ ,
    \new_Sorter100|12813_ , \new_Sorter100|12814_ , \new_Sorter100|12815_ ,
    \new_Sorter100|12816_ , \new_Sorter100|12817_ , \new_Sorter100|12818_ ,
    \new_Sorter100|12819_ , \new_Sorter100|12820_ , \new_Sorter100|12821_ ,
    \new_Sorter100|12822_ , \new_Sorter100|12823_ , \new_Sorter100|12824_ ,
    \new_Sorter100|12825_ , \new_Sorter100|12826_ , \new_Sorter100|12827_ ,
    \new_Sorter100|12828_ , \new_Sorter100|12829_ , \new_Sorter100|12830_ ,
    \new_Sorter100|12831_ , \new_Sorter100|12832_ , \new_Sorter100|12833_ ,
    \new_Sorter100|12834_ , \new_Sorter100|12835_ , \new_Sorter100|12836_ ,
    \new_Sorter100|12837_ , \new_Sorter100|12838_ , \new_Sorter100|12839_ ,
    \new_Sorter100|12840_ , \new_Sorter100|12841_ , \new_Sorter100|12842_ ,
    \new_Sorter100|12843_ , \new_Sorter100|12844_ , \new_Sorter100|12845_ ,
    \new_Sorter100|12846_ , \new_Sorter100|12847_ , \new_Sorter100|12848_ ,
    \new_Sorter100|12849_ , \new_Sorter100|12850_ , \new_Sorter100|12851_ ,
    \new_Sorter100|12852_ , \new_Sorter100|12853_ , \new_Sorter100|12854_ ,
    \new_Sorter100|12855_ , \new_Sorter100|12856_ , \new_Sorter100|12857_ ,
    \new_Sorter100|12858_ , \new_Sorter100|12859_ , \new_Sorter100|12860_ ,
    \new_Sorter100|12861_ , \new_Sorter100|12862_ , \new_Sorter100|12863_ ,
    \new_Sorter100|12864_ , \new_Sorter100|12865_ , \new_Sorter100|12866_ ,
    \new_Sorter100|12867_ , \new_Sorter100|12868_ , \new_Sorter100|12869_ ,
    \new_Sorter100|12870_ , \new_Sorter100|12871_ , \new_Sorter100|12872_ ,
    \new_Sorter100|12873_ , \new_Sorter100|12874_ , \new_Sorter100|12875_ ,
    \new_Sorter100|12876_ , \new_Sorter100|12877_ , \new_Sorter100|12878_ ,
    \new_Sorter100|12879_ , \new_Sorter100|12880_ , \new_Sorter100|12881_ ,
    \new_Sorter100|12882_ , \new_Sorter100|12883_ , \new_Sorter100|12884_ ,
    \new_Sorter100|12885_ , \new_Sorter100|12886_ , \new_Sorter100|12887_ ,
    \new_Sorter100|12888_ , \new_Sorter100|12889_ , \new_Sorter100|12890_ ,
    \new_Sorter100|12891_ , \new_Sorter100|12892_ , \new_Sorter100|12893_ ,
    \new_Sorter100|12894_ , \new_Sorter100|12895_ , \new_Sorter100|12896_ ,
    \new_Sorter100|12897_ , \new_Sorter100|12898_ , \new_Sorter100|12899_ ,
    \new_Sorter100|12900_ , \new_Sorter100|12999_ , \new_Sorter100|12901_ ,
    \new_Sorter100|12902_ , \new_Sorter100|12903_ , \new_Sorter100|12904_ ,
    \new_Sorter100|12905_ , \new_Sorter100|12906_ , \new_Sorter100|12907_ ,
    \new_Sorter100|12908_ , \new_Sorter100|12909_ , \new_Sorter100|12910_ ,
    \new_Sorter100|12911_ , \new_Sorter100|12912_ , \new_Sorter100|12913_ ,
    \new_Sorter100|12914_ , \new_Sorter100|12915_ , \new_Sorter100|12916_ ,
    \new_Sorter100|12917_ , \new_Sorter100|12918_ , \new_Sorter100|12919_ ,
    \new_Sorter100|12920_ , \new_Sorter100|12921_ , \new_Sorter100|12922_ ,
    \new_Sorter100|12923_ , \new_Sorter100|12924_ , \new_Sorter100|12925_ ,
    \new_Sorter100|12926_ , \new_Sorter100|12927_ , \new_Sorter100|12928_ ,
    \new_Sorter100|12929_ , \new_Sorter100|12930_ , \new_Sorter100|12931_ ,
    \new_Sorter100|12932_ , \new_Sorter100|12933_ , \new_Sorter100|12934_ ,
    \new_Sorter100|12935_ , \new_Sorter100|12936_ , \new_Sorter100|12937_ ,
    \new_Sorter100|12938_ , \new_Sorter100|12939_ , \new_Sorter100|12940_ ,
    \new_Sorter100|12941_ , \new_Sorter100|12942_ , \new_Sorter100|12943_ ,
    \new_Sorter100|12944_ , \new_Sorter100|12945_ , \new_Sorter100|12946_ ,
    \new_Sorter100|12947_ , \new_Sorter100|12948_ , \new_Sorter100|12949_ ,
    \new_Sorter100|12950_ , \new_Sorter100|12951_ , \new_Sorter100|12952_ ,
    \new_Sorter100|12953_ , \new_Sorter100|12954_ , \new_Sorter100|12955_ ,
    \new_Sorter100|12956_ , \new_Sorter100|12957_ , \new_Sorter100|12958_ ,
    \new_Sorter100|12959_ , \new_Sorter100|12960_ , \new_Sorter100|12961_ ,
    \new_Sorter100|12962_ , \new_Sorter100|12963_ , \new_Sorter100|12964_ ,
    \new_Sorter100|12965_ , \new_Sorter100|12966_ , \new_Sorter100|12967_ ,
    \new_Sorter100|12968_ , \new_Sorter100|12969_ , \new_Sorter100|12970_ ,
    \new_Sorter100|12971_ , \new_Sorter100|12972_ , \new_Sorter100|12973_ ,
    \new_Sorter100|12974_ , \new_Sorter100|12975_ , \new_Sorter100|12976_ ,
    \new_Sorter100|12977_ , \new_Sorter100|12978_ , \new_Sorter100|12979_ ,
    \new_Sorter100|12980_ , \new_Sorter100|12981_ , \new_Sorter100|12982_ ,
    \new_Sorter100|12983_ , \new_Sorter100|12984_ , \new_Sorter100|12985_ ,
    \new_Sorter100|12986_ , \new_Sorter100|12987_ , \new_Sorter100|12988_ ,
    \new_Sorter100|12989_ , \new_Sorter100|12990_ , \new_Sorter100|12991_ ,
    \new_Sorter100|12992_ , \new_Sorter100|12993_ , \new_Sorter100|12994_ ,
    \new_Sorter100|12995_ , \new_Sorter100|12996_ , \new_Sorter100|12997_ ,
    \new_Sorter100|12998_ , \new_Sorter100|13000_ , \new_Sorter100|13001_ ,
    \new_Sorter100|13002_ , \new_Sorter100|13003_ , \new_Sorter100|13004_ ,
    \new_Sorter100|13005_ , \new_Sorter100|13006_ , \new_Sorter100|13007_ ,
    \new_Sorter100|13008_ , \new_Sorter100|13009_ , \new_Sorter100|13010_ ,
    \new_Sorter100|13011_ , \new_Sorter100|13012_ , \new_Sorter100|13013_ ,
    \new_Sorter100|13014_ , \new_Sorter100|13015_ , \new_Sorter100|13016_ ,
    \new_Sorter100|13017_ , \new_Sorter100|13018_ , \new_Sorter100|13019_ ,
    \new_Sorter100|13020_ , \new_Sorter100|13021_ , \new_Sorter100|13022_ ,
    \new_Sorter100|13023_ , \new_Sorter100|13024_ , \new_Sorter100|13025_ ,
    \new_Sorter100|13026_ , \new_Sorter100|13027_ , \new_Sorter100|13028_ ,
    \new_Sorter100|13029_ , \new_Sorter100|13030_ , \new_Sorter100|13031_ ,
    \new_Sorter100|13032_ , \new_Sorter100|13033_ , \new_Sorter100|13034_ ,
    \new_Sorter100|13035_ , \new_Sorter100|13036_ , \new_Sorter100|13037_ ,
    \new_Sorter100|13038_ , \new_Sorter100|13039_ , \new_Sorter100|13040_ ,
    \new_Sorter100|13041_ , \new_Sorter100|13042_ , \new_Sorter100|13043_ ,
    \new_Sorter100|13044_ , \new_Sorter100|13045_ , \new_Sorter100|13046_ ,
    \new_Sorter100|13047_ , \new_Sorter100|13048_ , \new_Sorter100|13049_ ,
    \new_Sorter100|13050_ , \new_Sorter100|13051_ , \new_Sorter100|13052_ ,
    \new_Sorter100|13053_ , \new_Sorter100|13054_ , \new_Sorter100|13055_ ,
    \new_Sorter100|13056_ , \new_Sorter100|13057_ , \new_Sorter100|13058_ ,
    \new_Sorter100|13059_ , \new_Sorter100|13060_ , \new_Sorter100|13061_ ,
    \new_Sorter100|13062_ , \new_Sorter100|13063_ , \new_Sorter100|13064_ ,
    \new_Sorter100|13065_ , \new_Sorter100|13066_ , \new_Sorter100|13067_ ,
    \new_Sorter100|13068_ , \new_Sorter100|13069_ , \new_Sorter100|13070_ ,
    \new_Sorter100|13071_ , \new_Sorter100|13072_ , \new_Sorter100|13073_ ,
    \new_Sorter100|13074_ , \new_Sorter100|13075_ , \new_Sorter100|13076_ ,
    \new_Sorter100|13077_ , \new_Sorter100|13078_ , \new_Sorter100|13079_ ,
    \new_Sorter100|13080_ , \new_Sorter100|13081_ , \new_Sorter100|13082_ ,
    \new_Sorter100|13083_ , \new_Sorter100|13084_ , \new_Sorter100|13085_ ,
    \new_Sorter100|13086_ , \new_Sorter100|13087_ , \new_Sorter100|13088_ ,
    \new_Sorter100|13089_ , \new_Sorter100|13090_ , \new_Sorter100|13091_ ,
    \new_Sorter100|13092_ , \new_Sorter100|13093_ , \new_Sorter100|13094_ ,
    \new_Sorter100|13095_ , \new_Sorter100|13096_ , \new_Sorter100|13097_ ,
    \new_Sorter100|13098_ , \new_Sorter100|13099_ , \new_Sorter100|13100_ ,
    \new_Sorter100|13199_ , \new_Sorter100|13101_ , \new_Sorter100|13102_ ,
    \new_Sorter100|13103_ , \new_Sorter100|13104_ , \new_Sorter100|13105_ ,
    \new_Sorter100|13106_ , \new_Sorter100|13107_ , \new_Sorter100|13108_ ,
    \new_Sorter100|13109_ , \new_Sorter100|13110_ , \new_Sorter100|13111_ ,
    \new_Sorter100|13112_ , \new_Sorter100|13113_ , \new_Sorter100|13114_ ,
    \new_Sorter100|13115_ , \new_Sorter100|13116_ , \new_Sorter100|13117_ ,
    \new_Sorter100|13118_ , \new_Sorter100|13119_ , \new_Sorter100|13120_ ,
    \new_Sorter100|13121_ , \new_Sorter100|13122_ , \new_Sorter100|13123_ ,
    \new_Sorter100|13124_ , \new_Sorter100|13125_ , \new_Sorter100|13126_ ,
    \new_Sorter100|13127_ , \new_Sorter100|13128_ , \new_Sorter100|13129_ ,
    \new_Sorter100|13130_ , \new_Sorter100|13131_ , \new_Sorter100|13132_ ,
    \new_Sorter100|13133_ , \new_Sorter100|13134_ , \new_Sorter100|13135_ ,
    \new_Sorter100|13136_ , \new_Sorter100|13137_ , \new_Sorter100|13138_ ,
    \new_Sorter100|13139_ , \new_Sorter100|13140_ , \new_Sorter100|13141_ ,
    \new_Sorter100|13142_ , \new_Sorter100|13143_ , \new_Sorter100|13144_ ,
    \new_Sorter100|13145_ , \new_Sorter100|13146_ , \new_Sorter100|13147_ ,
    \new_Sorter100|13148_ , \new_Sorter100|13149_ , \new_Sorter100|13150_ ,
    \new_Sorter100|13151_ , \new_Sorter100|13152_ , \new_Sorter100|13153_ ,
    \new_Sorter100|13154_ , \new_Sorter100|13155_ , \new_Sorter100|13156_ ,
    \new_Sorter100|13157_ , \new_Sorter100|13158_ , \new_Sorter100|13159_ ,
    \new_Sorter100|13160_ , \new_Sorter100|13161_ , \new_Sorter100|13162_ ,
    \new_Sorter100|13163_ , \new_Sorter100|13164_ , \new_Sorter100|13165_ ,
    \new_Sorter100|13166_ , \new_Sorter100|13167_ , \new_Sorter100|13168_ ,
    \new_Sorter100|13169_ , \new_Sorter100|13170_ , \new_Sorter100|13171_ ,
    \new_Sorter100|13172_ , \new_Sorter100|13173_ , \new_Sorter100|13174_ ,
    \new_Sorter100|13175_ , \new_Sorter100|13176_ , \new_Sorter100|13177_ ,
    \new_Sorter100|13178_ , \new_Sorter100|13179_ , \new_Sorter100|13180_ ,
    \new_Sorter100|13181_ , \new_Sorter100|13182_ , \new_Sorter100|13183_ ,
    \new_Sorter100|13184_ , \new_Sorter100|13185_ , \new_Sorter100|13186_ ,
    \new_Sorter100|13187_ , \new_Sorter100|13188_ , \new_Sorter100|13189_ ,
    \new_Sorter100|13190_ , \new_Sorter100|13191_ , \new_Sorter100|13192_ ,
    \new_Sorter100|13193_ , \new_Sorter100|13194_ , \new_Sorter100|13195_ ,
    \new_Sorter100|13196_ , \new_Sorter100|13197_ , \new_Sorter100|13198_ ,
    \new_Sorter100|13200_ , \new_Sorter100|13201_ , \new_Sorter100|13202_ ,
    \new_Sorter100|13203_ , \new_Sorter100|13204_ , \new_Sorter100|13205_ ,
    \new_Sorter100|13206_ , \new_Sorter100|13207_ , \new_Sorter100|13208_ ,
    \new_Sorter100|13209_ , \new_Sorter100|13210_ , \new_Sorter100|13211_ ,
    \new_Sorter100|13212_ , \new_Sorter100|13213_ , \new_Sorter100|13214_ ,
    \new_Sorter100|13215_ , \new_Sorter100|13216_ , \new_Sorter100|13217_ ,
    \new_Sorter100|13218_ , \new_Sorter100|13219_ , \new_Sorter100|13220_ ,
    \new_Sorter100|13221_ , \new_Sorter100|13222_ , \new_Sorter100|13223_ ,
    \new_Sorter100|13224_ , \new_Sorter100|13225_ , \new_Sorter100|13226_ ,
    \new_Sorter100|13227_ , \new_Sorter100|13228_ , \new_Sorter100|13229_ ,
    \new_Sorter100|13230_ , \new_Sorter100|13231_ , \new_Sorter100|13232_ ,
    \new_Sorter100|13233_ , \new_Sorter100|13234_ , \new_Sorter100|13235_ ,
    \new_Sorter100|13236_ , \new_Sorter100|13237_ , \new_Sorter100|13238_ ,
    \new_Sorter100|13239_ , \new_Sorter100|13240_ , \new_Sorter100|13241_ ,
    \new_Sorter100|13242_ , \new_Sorter100|13243_ , \new_Sorter100|13244_ ,
    \new_Sorter100|13245_ , \new_Sorter100|13246_ , \new_Sorter100|13247_ ,
    \new_Sorter100|13248_ , \new_Sorter100|13249_ , \new_Sorter100|13250_ ,
    \new_Sorter100|13251_ , \new_Sorter100|13252_ , \new_Sorter100|13253_ ,
    \new_Sorter100|13254_ , \new_Sorter100|13255_ , \new_Sorter100|13256_ ,
    \new_Sorter100|13257_ , \new_Sorter100|13258_ , \new_Sorter100|13259_ ,
    \new_Sorter100|13260_ , \new_Sorter100|13261_ , \new_Sorter100|13262_ ,
    \new_Sorter100|13263_ , \new_Sorter100|13264_ , \new_Sorter100|13265_ ,
    \new_Sorter100|13266_ , \new_Sorter100|13267_ , \new_Sorter100|13268_ ,
    \new_Sorter100|13269_ , \new_Sorter100|13270_ , \new_Sorter100|13271_ ,
    \new_Sorter100|13272_ , \new_Sorter100|13273_ , \new_Sorter100|13274_ ,
    \new_Sorter100|13275_ , \new_Sorter100|13276_ , \new_Sorter100|13277_ ,
    \new_Sorter100|13278_ , \new_Sorter100|13279_ , \new_Sorter100|13280_ ,
    \new_Sorter100|13281_ , \new_Sorter100|13282_ , \new_Sorter100|13283_ ,
    \new_Sorter100|13284_ , \new_Sorter100|13285_ , \new_Sorter100|13286_ ,
    \new_Sorter100|13287_ , \new_Sorter100|13288_ , \new_Sorter100|13289_ ,
    \new_Sorter100|13290_ , \new_Sorter100|13291_ , \new_Sorter100|13292_ ,
    \new_Sorter100|13293_ , \new_Sorter100|13294_ , \new_Sorter100|13295_ ,
    \new_Sorter100|13296_ , \new_Sorter100|13297_ , \new_Sorter100|13298_ ,
    \new_Sorter100|13299_ , \new_Sorter100|13300_ , \new_Sorter100|13399_ ,
    \new_Sorter100|13301_ , \new_Sorter100|13302_ , \new_Sorter100|13303_ ,
    \new_Sorter100|13304_ , \new_Sorter100|13305_ , \new_Sorter100|13306_ ,
    \new_Sorter100|13307_ , \new_Sorter100|13308_ , \new_Sorter100|13309_ ,
    \new_Sorter100|13310_ , \new_Sorter100|13311_ , \new_Sorter100|13312_ ,
    \new_Sorter100|13313_ , \new_Sorter100|13314_ , \new_Sorter100|13315_ ,
    \new_Sorter100|13316_ , \new_Sorter100|13317_ , \new_Sorter100|13318_ ,
    \new_Sorter100|13319_ , \new_Sorter100|13320_ , \new_Sorter100|13321_ ,
    \new_Sorter100|13322_ , \new_Sorter100|13323_ , \new_Sorter100|13324_ ,
    \new_Sorter100|13325_ , \new_Sorter100|13326_ , \new_Sorter100|13327_ ,
    \new_Sorter100|13328_ , \new_Sorter100|13329_ , \new_Sorter100|13330_ ,
    \new_Sorter100|13331_ , \new_Sorter100|13332_ , \new_Sorter100|13333_ ,
    \new_Sorter100|13334_ , \new_Sorter100|13335_ , \new_Sorter100|13336_ ,
    \new_Sorter100|13337_ , \new_Sorter100|13338_ , \new_Sorter100|13339_ ,
    \new_Sorter100|13340_ , \new_Sorter100|13341_ , \new_Sorter100|13342_ ,
    \new_Sorter100|13343_ , \new_Sorter100|13344_ , \new_Sorter100|13345_ ,
    \new_Sorter100|13346_ , \new_Sorter100|13347_ , \new_Sorter100|13348_ ,
    \new_Sorter100|13349_ , \new_Sorter100|13350_ , \new_Sorter100|13351_ ,
    \new_Sorter100|13352_ , \new_Sorter100|13353_ , \new_Sorter100|13354_ ,
    \new_Sorter100|13355_ , \new_Sorter100|13356_ , \new_Sorter100|13357_ ,
    \new_Sorter100|13358_ , \new_Sorter100|13359_ , \new_Sorter100|13360_ ,
    \new_Sorter100|13361_ , \new_Sorter100|13362_ , \new_Sorter100|13363_ ,
    \new_Sorter100|13364_ , \new_Sorter100|13365_ , \new_Sorter100|13366_ ,
    \new_Sorter100|13367_ , \new_Sorter100|13368_ , \new_Sorter100|13369_ ,
    \new_Sorter100|13370_ , \new_Sorter100|13371_ , \new_Sorter100|13372_ ,
    \new_Sorter100|13373_ , \new_Sorter100|13374_ , \new_Sorter100|13375_ ,
    \new_Sorter100|13376_ , \new_Sorter100|13377_ , \new_Sorter100|13378_ ,
    \new_Sorter100|13379_ , \new_Sorter100|13380_ , \new_Sorter100|13381_ ,
    \new_Sorter100|13382_ , \new_Sorter100|13383_ , \new_Sorter100|13384_ ,
    \new_Sorter100|13385_ , \new_Sorter100|13386_ , \new_Sorter100|13387_ ,
    \new_Sorter100|13388_ , \new_Sorter100|13389_ , \new_Sorter100|13390_ ,
    \new_Sorter100|13391_ , \new_Sorter100|13392_ , \new_Sorter100|13393_ ,
    \new_Sorter100|13394_ , \new_Sorter100|13395_ , \new_Sorter100|13396_ ,
    \new_Sorter100|13397_ , \new_Sorter100|13398_ , \new_Sorter100|13400_ ,
    \new_Sorter100|13401_ , \new_Sorter100|13402_ , \new_Sorter100|13403_ ,
    \new_Sorter100|13404_ , \new_Sorter100|13405_ , \new_Sorter100|13406_ ,
    \new_Sorter100|13407_ , \new_Sorter100|13408_ , \new_Sorter100|13409_ ,
    \new_Sorter100|13410_ , \new_Sorter100|13411_ , \new_Sorter100|13412_ ,
    \new_Sorter100|13413_ , \new_Sorter100|13414_ , \new_Sorter100|13415_ ,
    \new_Sorter100|13416_ , \new_Sorter100|13417_ , \new_Sorter100|13418_ ,
    \new_Sorter100|13419_ , \new_Sorter100|13420_ , \new_Sorter100|13421_ ,
    \new_Sorter100|13422_ , \new_Sorter100|13423_ , \new_Sorter100|13424_ ,
    \new_Sorter100|13425_ , \new_Sorter100|13426_ , \new_Sorter100|13427_ ,
    \new_Sorter100|13428_ , \new_Sorter100|13429_ , \new_Sorter100|13430_ ,
    \new_Sorter100|13431_ , \new_Sorter100|13432_ , \new_Sorter100|13433_ ,
    \new_Sorter100|13434_ , \new_Sorter100|13435_ , \new_Sorter100|13436_ ,
    \new_Sorter100|13437_ , \new_Sorter100|13438_ , \new_Sorter100|13439_ ,
    \new_Sorter100|13440_ , \new_Sorter100|13441_ , \new_Sorter100|13442_ ,
    \new_Sorter100|13443_ , \new_Sorter100|13444_ , \new_Sorter100|13445_ ,
    \new_Sorter100|13446_ , \new_Sorter100|13447_ , \new_Sorter100|13448_ ,
    \new_Sorter100|13449_ , \new_Sorter100|13450_ , \new_Sorter100|13451_ ,
    \new_Sorter100|13452_ , \new_Sorter100|13453_ , \new_Sorter100|13454_ ,
    \new_Sorter100|13455_ , \new_Sorter100|13456_ , \new_Sorter100|13457_ ,
    \new_Sorter100|13458_ , \new_Sorter100|13459_ , \new_Sorter100|13460_ ,
    \new_Sorter100|13461_ , \new_Sorter100|13462_ , \new_Sorter100|13463_ ,
    \new_Sorter100|13464_ , \new_Sorter100|13465_ , \new_Sorter100|13466_ ,
    \new_Sorter100|13467_ , \new_Sorter100|13468_ , \new_Sorter100|13469_ ,
    \new_Sorter100|13470_ , \new_Sorter100|13471_ , \new_Sorter100|13472_ ,
    \new_Sorter100|13473_ , \new_Sorter100|13474_ , \new_Sorter100|13475_ ,
    \new_Sorter100|13476_ , \new_Sorter100|13477_ , \new_Sorter100|13478_ ,
    \new_Sorter100|13479_ , \new_Sorter100|13480_ , \new_Sorter100|13481_ ,
    \new_Sorter100|13482_ , \new_Sorter100|13483_ , \new_Sorter100|13484_ ,
    \new_Sorter100|13485_ , \new_Sorter100|13486_ , \new_Sorter100|13487_ ,
    \new_Sorter100|13488_ , \new_Sorter100|13489_ , \new_Sorter100|13490_ ,
    \new_Sorter100|13491_ , \new_Sorter100|13492_ , \new_Sorter100|13493_ ,
    \new_Sorter100|13494_ , \new_Sorter100|13495_ , \new_Sorter100|13496_ ,
    \new_Sorter100|13497_ , \new_Sorter100|13498_ , \new_Sorter100|13499_ ,
    \new_Sorter100|13500_ , \new_Sorter100|13599_ , \new_Sorter100|13501_ ,
    \new_Sorter100|13502_ , \new_Sorter100|13503_ , \new_Sorter100|13504_ ,
    \new_Sorter100|13505_ , \new_Sorter100|13506_ , \new_Sorter100|13507_ ,
    \new_Sorter100|13508_ , \new_Sorter100|13509_ , \new_Sorter100|13510_ ,
    \new_Sorter100|13511_ , \new_Sorter100|13512_ , \new_Sorter100|13513_ ,
    \new_Sorter100|13514_ , \new_Sorter100|13515_ , \new_Sorter100|13516_ ,
    \new_Sorter100|13517_ , \new_Sorter100|13518_ , \new_Sorter100|13519_ ,
    \new_Sorter100|13520_ , \new_Sorter100|13521_ , \new_Sorter100|13522_ ,
    \new_Sorter100|13523_ , \new_Sorter100|13524_ , \new_Sorter100|13525_ ,
    \new_Sorter100|13526_ , \new_Sorter100|13527_ , \new_Sorter100|13528_ ,
    \new_Sorter100|13529_ , \new_Sorter100|13530_ , \new_Sorter100|13531_ ,
    \new_Sorter100|13532_ , \new_Sorter100|13533_ , \new_Sorter100|13534_ ,
    \new_Sorter100|13535_ , \new_Sorter100|13536_ , \new_Sorter100|13537_ ,
    \new_Sorter100|13538_ , \new_Sorter100|13539_ , \new_Sorter100|13540_ ,
    \new_Sorter100|13541_ , \new_Sorter100|13542_ , \new_Sorter100|13543_ ,
    \new_Sorter100|13544_ , \new_Sorter100|13545_ , \new_Sorter100|13546_ ,
    \new_Sorter100|13547_ , \new_Sorter100|13548_ , \new_Sorter100|13549_ ,
    \new_Sorter100|13550_ , \new_Sorter100|13551_ , \new_Sorter100|13552_ ,
    \new_Sorter100|13553_ , \new_Sorter100|13554_ , \new_Sorter100|13555_ ,
    \new_Sorter100|13556_ , \new_Sorter100|13557_ , \new_Sorter100|13558_ ,
    \new_Sorter100|13559_ , \new_Sorter100|13560_ , \new_Sorter100|13561_ ,
    \new_Sorter100|13562_ , \new_Sorter100|13563_ , \new_Sorter100|13564_ ,
    \new_Sorter100|13565_ , \new_Sorter100|13566_ , \new_Sorter100|13567_ ,
    \new_Sorter100|13568_ , \new_Sorter100|13569_ , \new_Sorter100|13570_ ,
    \new_Sorter100|13571_ , \new_Sorter100|13572_ , \new_Sorter100|13573_ ,
    \new_Sorter100|13574_ , \new_Sorter100|13575_ , \new_Sorter100|13576_ ,
    \new_Sorter100|13577_ , \new_Sorter100|13578_ , \new_Sorter100|13579_ ,
    \new_Sorter100|13580_ , \new_Sorter100|13581_ , \new_Sorter100|13582_ ,
    \new_Sorter100|13583_ , \new_Sorter100|13584_ , \new_Sorter100|13585_ ,
    \new_Sorter100|13586_ , \new_Sorter100|13587_ , \new_Sorter100|13588_ ,
    \new_Sorter100|13589_ , \new_Sorter100|13590_ , \new_Sorter100|13591_ ,
    \new_Sorter100|13592_ , \new_Sorter100|13593_ , \new_Sorter100|13594_ ,
    \new_Sorter100|13595_ , \new_Sorter100|13596_ , \new_Sorter100|13597_ ,
    \new_Sorter100|13598_ , \new_Sorter100|13600_ , \new_Sorter100|13601_ ,
    \new_Sorter100|13602_ , \new_Sorter100|13603_ , \new_Sorter100|13604_ ,
    \new_Sorter100|13605_ , \new_Sorter100|13606_ , \new_Sorter100|13607_ ,
    \new_Sorter100|13608_ , \new_Sorter100|13609_ , \new_Sorter100|13610_ ,
    \new_Sorter100|13611_ , \new_Sorter100|13612_ , \new_Sorter100|13613_ ,
    \new_Sorter100|13614_ , \new_Sorter100|13615_ , \new_Sorter100|13616_ ,
    \new_Sorter100|13617_ , \new_Sorter100|13618_ , \new_Sorter100|13619_ ,
    \new_Sorter100|13620_ , \new_Sorter100|13621_ , \new_Sorter100|13622_ ,
    \new_Sorter100|13623_ , \new_Sorter100|13624_ , \new_Sorter100|13625_ ,
    \new_Sorter100|13626_ , \new_Sorter100|13627_ , \new_Sorter100|13628_ ,
    \new_Sorter100|13629_ , \new_Sorter100|13630_ , \new_Sorter100|13631_ ,
    \new_Sorter100|13632_ , \new_Sorter100|13633_ , \new_Sorter100|13634_ ,
    \new_Sorter100|13635_ , \new_Sorter100|13636_ , \new_Sorter100|13637_ ,
    \new_Sorter100|13638_ , \new_Sorter100|13639_ , \new_Sorter100|13640_ ,
    \new_Sorter100|13641_ , \new_Sorter100|13642_ , \new_Sorter100|13643_ ,
    \new_Sorter100|13644_ , \new_Sorter100|13645_ , \new_Sorter100|13646_ ,
    \new_Sorter100|13647_ , \new_Sorter100|13648_ , \new_Sorter100|13649_ ,
    \new_Sorter100|13650_ , \new_Sorter100|13651_ , \new_Sorter100|13652_ ,
    \new_Sorter100|13653_ , \new_Sorter100|13654_ , \new_Sorter100|13655_ ,
    \new_Sorter100|13656_ , \new_Sorter100|13657_ , \new_Sorter100|13658_ ,
    \new_Sorter100|13659_ , \new_Sorter100|13660_ , \new_Sorter100|13661_ ,
    \new_Sorter100|13662_ , \new_Sorter100|13663_ , \new_Sorter100|13664_ ,
    \new_Sorter100|13665_ , \new_Sorter100|13666_ , \new_Sorter100|13667_ ,
    \new_Sorter100|13668_ , \new_Sorter100|13669_ , \new_Sorter100|13670_ ,
    \new_Sorter100|13671_ , \new_Sorter100|13672_ , \new_Sorter100|13673_ ,
    \new_Sorter100|13674_ , \new_Sorter100|13675_ , \new_Sorter100|13676_ ,
    \new_Sorter100|13677_ , \new_Sorter100|13678_ , \new_Sorter100|13679_ ,
    \new_Sorter100|13680_ , \new_Sorter100|13681_ , \new_Sorter100|13682_ ,
    \new_Sorter100|13683_ , \new_Sorter100|13684_ , \new_Sorter100|13685_ ,
    \new_Sorter100|13686_ , \new_Sorter100|13687_ , \new_Sorter100|13688_ ,
    \new_Sorter100|13689_ , \new_Sorter100|13690_ , \new_Sorter100|13691_ ,
    \new_Sorter100|13692_ , \new_Sorter100|13693_ , \new_Sorter100|13694_ ,
    \new_Sorter100|13695_ , \new_Sorter100|13696_ , \new_Sorter100|13697_ ,
    \new_Sorter100|13698_ , \new_Sorter100|13699_ , \new_Sorter100|13700_ ,
    \new_Sorter100|13799_ , \new_Sorter100|13701_ , \new_Sorter100|13702_ ,
    \new_Sorter100|13703_ , \new_Sorter100|13704_ , \new_Sorter100|13705_ ,
    \new_Sorter100|13706_ , \new_Sorter100|13707_ , \new_Sorter100|13708_ ,
    \new_Sorter100|13709_ , \new_Sorter100|13710_ , \new_Sorter100|13711_ ,
    \new_Sorter100|13712_ , \new_Sorter100|13713_ , \new_Sorter100|13714_ ,
    \new_Sorter100|13715_ , \new_Sorter100|13716_ , \new_Sorter100|13717_ ,
    \new_Sorter100|13718_ , \new_Sorter100|13719_ , \new_Sorter100|13720_ ,
    \new_Sorter100|13721_ , \new_Sorter100|13722_ , \new_Sorter100|13723_ ,
    \new_Sorter100|13724_ , \new_Sorter100|13725_ , \new_Sorter100|13726_ ,
    \new_Sorter100|13727_ , \new_Sorter100|13728_ , \new_Sorter100|13729_ ,
    \new_Sorter100|13730_ , \new_Sorter100|13731_ , \new_Sorter100|13732_ ,
    \new_Sorter100|13733_ , \new_Sorter100|13734_ , \new_Sorter100|13735_ ,
    \new_Sorter100|13736_ , \new_Sorter100|13737_ , \new_Sorter100|13738_ ,
    \new_Sorter100|13739_ , \new_Sorter100|13740_ , \new_Sorter100|13741_ ,
    \new_Sorter100|13742_ , \new_Sorter100|13743_ , \new_Sorter100|13744_ ,
    \new_Sorter100|13745_ , \new_Sorter100|13746_ , \new_Sorter100|13747_ ,
    \new_Sorter100|13748_ , \new_Sorter100|13749_ , \new_Sorter100|13750_ ,
    \new_Sorter100|13751_ , \new_Sorter100|13752_ , \new_Sorter100|13753_ ,
    \new_Sorter100|13754_ , \new_Sorter100|13755_ , \new_Sorter100|13756_ ,
    \new_Sorter100|13757_ , \new_Sorter100|13758_ , \new_Sorter100|13759_ ,
    \new_Sorter100|13760_ , \new_Sorter100|13761_ , \new_Sorter100|13762_ ,
    \new_Sorter100|13763_ , \new_Sorter100|13764_ , \new_Sorter100|13765_ ,
    \new_Sorter100|13766_ , \new_Sorter100|13767_ , \new_Sorter100|13768_ ,
    \new_Sorter100|13769_ , \new_Sorter100|13770_ , \new_Sorter100|13771_ ,
    \new_Sorter100|13772_ , \new_Sorter100|13773_ , \new_Sorter100|13774_ ,
    \new_Sorter100|13775_ , \new_Sorter100|13776_ , \new_Sorter100|13777_ ,
    \new_Sorter100|13778_ , \new_Sorter100|13779_ , \new_Sorter100|13780_ ,
    \new_Sorter100|13781_ , \new_Sorter100|13782_ , \new_Sorter100|13783_ ,
    \new_Sorter100|13784_ , \new_Sorter100|13785_ , \new_Sorter100|13786_ ,
    \new_Sorter100|13787_ , \new_Sorter100|13788_ , \new_Sorter100|13789_ ,
    \new_Sorter100|13790_ , \new_Sorter100|13791_ , \new_Sorter100|13792_ ,
    \new_Sorter100|13793_ , \new_Sorter100|13794_ , \new_Sorter100|13795_ ,
    \new_Sorter100|13796_ , \new_Sorter100|13797_ , \new_Sorter100|13798_ ,
    \new_Sorter100|13800_ , \new_Sorter100|13801_ , \new_Sorter100|13802_ ,
    \new_Sorter100|13803_ , \new_Sorter100|13804_ , \new_Sorter100|13805_ ,
    \new_Sorter100|13806_ , \new_Sorter100|13807_ , \new_Sorter100|13808_ ,
    \new_Sorter100|13809_ , \new_Sorter100|13810_ , \new_Sorter100|13811_ ,
    \new_Sorter100|13812_ , \new_Sorter100|13813_ , \new_Sorter100|13814_ ,
    \new_Sorter100|13815_ , \new_Sorter100|13816_ , \new_Sorter100|13817_ ,
    \new_Sorter100|13818_ , \new_Sorter100|13819_ , \new_Sorter100|13820_ ,
    \new_Sorter100|13821_ , \new_Sorter100|13822_ , \new_Sorter100|13823_ ,
    \new_Sorter100|13824_ , \new_Sorter100|13825_ , \new_Sorter100|13826_ ,
    \new_Sorter100|13827_ , \new_Sorter100|13828_ , \new_Sorter100|13829_ ,
    \new_Sorter100|13830_ , \new_Sorter100|13831_ , \new_Sorter100|13832_ ,
    \new_Sorter100|13833_ , \new_Sorter100|13834_ , \new_Sorter100|13835_ ,
    \new_Sorter100|13836_ , \new_Sorter100|13837_ , \new_Sorter100|13838_ ,
    \new_Sorter100|13839_ , \new_Sorter100|13840_ , \new_Sorter100|13841_ ,
    \new_Sorter100|13842_ , \new_Sorter100|13843_ , \new_Sorter100|13844_ ,
    \new_Sorter100|13845_ , \new_Sorter100|13846_ , \new_Sorter100|13847_ ,
    \new_Sorter100|13848_ , \new_Sorter100|13849_ , \new_Sorter100|13850_ ,
    \new_Sorter100|13851_ , \new_Sorter100|13852_ , \new_Sorter100|13853_ ,
    \new_Sorter100|13854_ , \new_Sorter100|13855_ , \new_Sorter100|13856_ ,
    \new_Sorter100|13857_ , \new_Sorter100|13858_ , \new_Sorter100|13859_ ,
    \new_Sorter100|13860_ , \new_Sorter100|13861_ , \new_Sorter100|13862_ ,
    \new_Sorter100|13863_ , \new_Sorter100|13864_ , \new_Sorter100|13865_ ,
    \new_Sorter100|13866_ , \new_Sorter100|13867_ , \new_Sorter100|13868_ ,
    \new_Sorter100|13869_ , \new_Sorter100|13870_ , \new_Sorter100|13871_ ,
    \new_Sorter100|13872_ , \new_Sorter100|13873_ , \new_Sorter100|13874_ ,
    \new_Sorter100|13875_ , \new_Sorter100|13876_ , \new_Sorter100|13877_ ,
    \new_Sorter100|13878_ , \new_Sorter100|13879_ , \new_Sorter100|13880_ ,
    \new_Sorter100|13881_ , \new_Sorter100|13882_ , \new_Sorter100|13883_ ,
    \new_Sorter100|13884_ , \new_Sorter100|13885_ , \new_Sorter100|13886_ ,
    \new_Sorter100|13887_ , \new_Sorter100|13888_ , \new_Sorter100|13889_ ,
    \new_Sorter100|13890_ , \new_Sorter100|13891_ , \new_Sorter100|13892_ ,
    \new_Sorter100|13893_ , \new_Sorter100|13894_ , \new_Sorter100|13895_ ,
    \new_Sorter100|13896_ , \new_Sorter100|13897_ , \new_Sorter100|13898_ ,
    \new_Sorter100|13899_ , \new_Sorter100|13900_ , \new_Sorter100|13999_ ,
    \new_Sorter100|13901_ , \new_Sorter100|13902_ , \new_Sorter100|13903_ ,
    \new_Sorter100|13904_ , \new_Sorter100|13905_ , \new_Sorter100|13906_ ,
    \new_Sorter100|13907_ , \new_Sorter100|13908_ , \new_Sorter100|13909_ ,
    \new_Sorter100|13910_ , \new_Sorter100|13911_ , \new_Sorter100|13912_ ,
    \new_Sorter100|13913_ , \new_Sorter100|13914_ , \new_Sorter100|13915_ ,
    \new_Sorter100|13916_ , \new_Sorter100|13917_ , \new_Sorter100|13918_ ,
    \new_Sorter100|13919_ , \new_Sorter100|13920_ , \new_Sorter100|13921_ ,
    \new_Sorter100|13922_ , \new_Sorter100|13923_ , \new_Sorter100|13924_ ,
    \new_Sorter100|13925_ , \new_Sorter100|13926_ , \new_Sorter100|13927_ ,
    \new_Sorter100|13928_ , \new_Sorter100|13929_ , \new_Sorter100|13930_ ,
    \new_Sorter100|13931_ , \new_Sorter100|13932_ , \new_Sorter100|13933_ ,
    \new_Sorter100|13934_ , \new_Sorter100|13935_ , \new_Sorter100|13936_ ,
    \new_Sorter100|13937_ , \new_Sorter100|13938_ , \new_Sorter100|13939_ ,
    \new_Sorter100|13940_ , \new_Sorter100|13941_ , \new_Sorter100|13942_ ,
    \new_Sorter100|13943_ , \new_Sorter100|13944_ , \new_Sorter100|13945_ ,
    \new_Sorter100|13946_ , \new_Sorter100|13947_ , \new_Sorter100|13948_ ,
    \new_Sorter100|13949_ , \new_Sorter100|13950_ , \new_Sorter100|13951_ ,
    \new_Sorter100|13952_ , \new_Sorter100|13953_ , \new_Sorter100|13954_ ,
    \new_Sorter100|13955_ , \new_Sorter100|13956_ , \new_Sorter100|13957_ ,
    \new_Sorter100|13958_ , \new_Sorter100|13959_ , \new_Sorter100|13960_ ,
    \new_Sorter100|13961_ , \new_Sorter100|13962_ , \new_Sorter100|13963_ ,
    \new_Sorter100|13964_ , \new_Sorter100|13965_ , \new_Sorter100|13966_ ,
    \new_Sorter100|13967_ , \new_Sorter100|13968_ , \new_Sorter100|13969_ ,
    \new_Sorter100|13970_ , \new_Sorter100|13971_ , \new_Sorter100|13972_ ,
    \new_Sorter100|13973_ , \new_Sorter100|13974_ , \new_Sorter100|13975_ ,
    \new_Sorter100|13976_ , \new_Sorter100|13977_ , \new_Sorter100|13978_ ,
    \new_Sorter100|13979_ , \new_Sorter100|13980_ , \new_Sorter100|13981_ ,
    \new_Sorter100|13982_ , \new_Sorter100|13983_ , \new_Sorter100|13984_ ,
    \new_Sorter100|13985_ , \new_Sorter100|13986_ , \new_Sorter100|13987_ ,
    \new_Sorter100|13988_ , \new_Sorter100|13989_ , \new_Sorter100|13990_ ,
    \new_Sorter100|13991_ , \new_Sorter100|13992_ , \new_Sorter100|13993_ ,
    \new_Sorter100|13994_ , \new_Sorter100|13995_ , \new_Sorter100|13996_ ,
    \new_Sorter100|13997_ , \new_Sorter100|13998_ , \new_Sorter100|14000_ ,
    \new_Sorter100|14001_ , \new_Sorter100|14002_ , \new_Sorter100|14003_ ,
    \new_Sorter100|14004_ , \new_Sorter100|14005_ , \new_Sorter100|14006_ ,
    \new_Sorter100|14007_ , \new_Sorter100|14008_ , \new_Sorter100|14009_ ,
    \new_Sorter100|14010_ , \new_Sorter100|14011_ , \new_Sorter100|14012_ ,
    \new_Sorter100|14013_ , \new_Sorter100|14014_ , \new_Sorter100|14015_ ,
    \new_Sorter100|14016_ , \new_Sorter100|14017_ , \new_Sorter100|14018_ ,
    \new_Sorter100|14019_ , \new_Sorter100|14020_ , \new_Sorter100|14021_ ,
    \new_Sorter100|14022_ , \new_Sorter100|14023_ , \new_Sorter100|14024_ ,
    \new_Sorter100|14025_ , \new_Sorter100|14026_ , \new_Sorter100|14027_ ,
    \new_Sorter100|14028_ , \new_Sorter100|14029_ , \new_Sorter100|14030_ ,
    \new_Sorter100|14031_ , \new_Sorter100|14032_ , \new_Sorter100|14033_ ,
    \new_Sorter100|14034_ , \new_Sorter100|14035_ , \new_Sorter100|14036_ ,
    \new_Sorter100|14037_ , \new_Sorter100|14038_ , \new_Sorter100|14039_ ,
    \new_Sorter100|14040_ , \new_Sorter100|14041_ , \new_Sorter100|14042_ ,
    \new_Sorter100|14043_ , \new_Sorter100|14044_ , \new_Sorter100|14045_ ,
    \new_Sorter100|14046_ , \new_Sorter100|14047_ , \new_Sorter100|14048_ ,
    \new_Sorter100|14049_ , \new_Sorter100|14050_ , \new_Sorter100|14051_ ,
    \new_Sorter100|14052_ , \new_Sorter100|14053_ , \new_Sorter100|14054_ ,
    \new_Sorter100|14055_ , \new_Sorter100|14056_ , \new_Sorter100|14057_ ,
    \new_Sorter100|14058_ , \new_Sorter100|14059_ , \new_Sorter100|14060_ ,
    \new_Sorter100|14061_ , \new_Sorter100|14062_ , \new_Sorter100|14063_ ,
    \new_Sorter100|14064_ , \new_Sorter100|14065_ , \new_Sorter100|14066_ ,
    \new_Sorter100|14067_ , \new_Sorter100|14068_ , \new_Sorter100|14069_ ,
    \new_Sorter100|14070_ , \new_Sorter100|14071_ , \new_Sorter100|14072_ ,
    \new_Sorter100|14073_ , \new_Sorter100|14074_ , \new_Sorter100|14075_ ,
    \new_Sorter100|14076_ , \new_Sorter100|14077_ , \new_Sorter100|14078_ ,
    \new_Sorter100|14079_ , \new_Sorter100|14080_ , \new_Sorter100|14081_ ,
    \new_Sorter100|14082_ , \new_Sorter100|14083_ , \new_Sorter100|14084_ ,
    \new_Sorter100|14085_ , \new_Sorter100|14086_ , \new_Sorter100|14087_ ,
    \new_Sorter100|14088_ , \new_Sorter100|14089_ , \new_Sorter100|14090_ ,
    \new_Sorter100|14091_ , \new_Sorter100|14092_ , \new_Sorter100|14093_ ,
    \new_Sorter100|14094_ , \new_Sorter100|14095_ , \new_Sorter100|14096_ ,
    \new_Sorter100|14097_ , \new_Sorter100|14098_ , \new_Sorter100|14099_ ,
    \new_Sorter100|14100_ , \new_Sorter100|14199_ , \new_Sorter100|14101_ ,
    \new_Sorter100|14102_ , \new_Sorter100|14103_ , \new_Sorter100|14104_ ,
    \new_Sorter100|14105_ , \new_Sorter100|14106_ , \new_Sorter100|14107_ ,
    \new_Sorter100|14108_ , \new_Sorter100|14109_ , \new_Sorter100|14110_ ,
    \new_Sorter100|14111_ , \new_Sorter100|14112_ , \new_Sorter100|14113_ ,
    \new_Sorter100|14114_ , \new_Sorter100|14115_ , \new_Sorter100|14116_ ,
    \new_Sorter100|14117_ , \new_Sorter100|14118_ , \new_Sorter100|14119_ ,
    \new_Sorter100|14120_ , \new_Sorter100|14121_ , \new_Sorter100|14122_ ,
    \new_Sorter100|14123_ , \new_Sorter100|14124_ , \new_Sorter100|14125_ ,
    \new_Sorter100|14126_ , \new_Sorter100|14127_ , \new_Sorter100|14128_ ,
    \new_Sorter100|14129_ , \new_Sorter100|14130_ , \new_Sorter100|14131_ ,
    \new_Sorter100|14132_ , \new_Sorter100|14133_ , \new_Sorter100|14134_ ,
    \new_Sorter100|14135_ , \new_Sorter100|14136_ , \new_Sorter100|14137_ ,
    \new_Sorter100|14138_ , \new_Sorter100|14139_ , \new_Sorter100|14140_ ,
    \new_Sorter100|14141_ , \new_Sorter100|14142_ , \new_Sorter100|14143_ ,
    \new_Sorter100|14144_ , \new_Sorter100|14145_ , \new_Sorter100|14146_ ,
    \new_Sorter100|14147_ , \new_Sorter100|14148_ , \new_Sorter100|14149_ ,
    \new_Sorter100|14150_ , \new_Sorter100|14151_ , \new_Sorter100|14152_ ,
    \new_Sorter100|14153_ , \new_Sorter100|14154_ , \new_Sorter100|14155_ ,
    \new_Sorter100|14156_ , \new_Sorter100|14157_ , \new_Sorter100|14158_ ,
    \new_Sorter100|14159_ , \new_Sorter100|14160_ , \new_Sorter100|14161_ ,
    \new_Sorter100|14162_ , \new_Sorter100|14163_ , \new_Sorter100|14164_ ,
    \new_Sorter100|14165_ , \new_Sorter100|14166_ , \new_Sorter100|14167_ ,
    \new_Sorter100|14168_ , \new_Sorter100|14169_ , \new_Sorter100|14170_ ,
    \new_Sorter100|14171_ , \new_Sorter100|14172_ , \new_Sorter100|14173_ ,
    \new_Sorter100|14174_ , \new_Sorter100|14175_ , \new_Sorter100|14176_ ,
    \new_Sorter100|14177_ , \new_Sorter100|14178_ , \new_Sorter100|14179_ ,
    \new_Sorter100|14180_ , \new_Sorter100|14181_ , \new_Sorter100|14182_ ,
    \new_Sorter100|14183_ , \new_Sorter100|14184_ , \new_Sorter100|14185_ ,
    \new_Sorter100|14186_ , \new_Sorter100|14187_ , \new_Sorter100|14188_ ,
    \new_Sorter100|14189_ , \new_Sorter100|14190_ , \new_Sorter100|14191_ ,
    \new_Sorter100|14192_ , \new_Sorter100|14193_ , \new_Sorter100|14194_ ,
    \new_Sorter100|14195_ , \new_Sorter100|14196_ , \new_Sorter100|14197_ ,
    \new_Sorter100|14198_ , \new_Sorter100|14200_ , \new_Sorter100|14201_ ,
    \new_Sorter100|14202_ , \new_Sorter100|14203_ , \new_Sorter100|14204_ ,
    \new_Sorter100|14205_ , \new_Sorter100|14206_ , \new_Sorter100|14207_ ,
    \new_Sorter100|14208_ , \new_Sorter100|14209_ , \new_Sorter100|14210_ ,
    \new_Sorter100|14211_ , \new_Sorter100|14212_ , \new_Sorter100|14213_ ,
    \new_Sorter100|14214_ , \new_Sorter100|14215_ , \new_Sorter100|14216_ ,
    \new_Sorter100|14217_ , \new_Sorter100|14218_ , \new_Sorter100|14219_ ,
    \new_Sorter100|14220_ , \new_Sorter100|14221_ , \new_Sorter100|14222_ ,
    \new_Sorter100|14223_ , \new_Sorter100|14224_ , \new_Sorter100|14225_ ,
    \new_Sorter100|14226_ , \new_Sorter100|14227_ , \new_Sorter100|14228_ ,
    \new_Sorter100|14229_ , \new_Sorter100|14230_ , \new_Sorter100|14231_ ,
    \new_Sorter100|14232_ , \new_Sorter100|14233_ , \new_Sorter100|14234_ ,
    \new_Sorter100|14235_ , \new_Sorter100|14236_ , \new_Sorter100|14237_ ,
    \new_Sorter100|14238_ , \new_Sorter100|14239_ , \new_Sorter100|14240_ ,
    \new_Sorter100|14241_ , \new_Sorter100|14242_ , \new_Sorter100|14243_ ,
    \new_Sorter100|14244_ , \new_Sorter100|14245_ , \new_Sorter100|14246_ ,
    \new_Sorter100|14247_ , \new_Sorter100|14248_ , \new_Sorter100|14249_ ,
    \new_Sorter100|14250_ , \new_Sorter100|14251_ , \new_Sorter100|14252_ ,
    \new_Sorter100|14253_ , \new_Sorter100|14254_ , \new_Sorter100|14255_ ,
    \new_Sorter100|14256_ , \new_Sorter100|14257_ , \new_Sorter100|14258_ ,
    \new_Sorter100|14259_ , \new_Sorter100|14260_ , \new_Sorter100|14261_ ,
    \new_Sorter100|14262_ , \new_Sorter100|14263_ , \new_Sorter100|14264_ ,
    \new_Sorter100|14265_ , \new_Sorter100|14266_ , \new_Sorter100|14267_ ,
    \new_Sorter100|14268_ , \new_Sorter100|14269_ , \new_Sorter100|14270_ ,
    \new_Sorter100|14271_ , \new_Sorter100|14272_ , \new_Sorter100|14273_ ,
    \new_Sorter100|14274_ , \new_Sorter100|14275_ , \new_Sorter100|14276_ ,
    \new_Sorter100|14277_ , \new_Sorter100|14278_ , \new_Sorter100|14279_ ,
    \new_Sorter100|14280_ , \new_Sorter100|14281_ , \new_Sorter100|14282_ ,
    \new_Sorter100|14283_ , \new_Sorter100|14284_ , \new_Sorter100|14285_ ,
    \new_Sorter100|14286_ , \new_Sorter100|14287_ , \new_Sorter100|14288_ ,
    \new_Sorter100|14289_ , \new_Sorter100|14290_ , \new_Sorter100|14291_ ,
    \new_Sorter100|14292_ , \new_Sorter100|14293_ , \new_Sorter100|14294_ ,
    \new_Sorter100|14295_ , \new_Sorter100|14296_ , \new_Sorter100|14297_ ,
    \new_Sorter100|14298_ , \new_Sorter100|14299_ , \new_Sorter100|14300_ ,
    \new_Sorter100|14399_ , \new_Sorter100|14301_ , \new_Sorter100|14302_ ,
    \new_Sorter100|14303_ , \new_Sorter100|14304_ , \new_Sorter100|14305_ ,
    \new_Sorter100|14306_ , \new_Sorter100|14307_ , \new_Sorter100|14308_ ,
    \new_Sorter100|14309_ , \new_Sorter100|14310_ , \new_Sorter100|14311_ ,
    \new_Sorter100|14312_ , \new_Sorter100|14313_ , \new_Sorter100|14314_ ,
    \new_Sorter100|14315_ , \new_Sorter100|14316_ , \new_Sorter100|14317_ ,
    \new_Sorter100|14318_ , \new_Sorter100|14319_ , \new_Sorter100|14320_ ,
    \new_Sorter100|14321_ , \new_Sorter100|14322_ , \new_Sorter100|14323_ ,
    \new_Sorter100|14324_ , \new_Sorter100|14325_ , \new_Sorter100|14326_ ,
    \new_Sorter100|14327_ , \new_Sorter100|14328_ , \new_Sorter100|14329_ ,
    \new_Sorter100|14330_ , \new_Sorter100|14331_ , \new_Sorter100|14332_ ,
    \new_Sorter100|14333_ , \new_Sorter100|14334_ , \new_Sorter100|14335_ ,
    \new_Sorter100|14336_ , \new_Sorter100|14337_ , \new_Sorter100|14338_ ,
    \new_Sorter100|14339_ , \new_Sorter100|14340_ , \new_Sorter100|14341_ ,
    \new_Sorter100|14342_ , \new_Sorter100|14343_ , \new_Sorter100|14344_ ,
    \new_Sorter100|14345_ , \new_Sorter100|14346_ , \new_Sorter100|14347_ ,
    \new_Sorter100|14348_ , \new_Sorter100|14349_ , \new_Sorter100|14350_ ,
    \new_Sorter100|14351_ , \new_Sorter100|14352_ , \new_Sorter100|14353_ ,
    \new_Sorter100|14354_ , \new_Sorter100|14355_ , \new_Sorter100|14356_ ,
    \new_Sorter100|14357_ , \new_Sorter100|14358_ , \new_Sorter100|14359_ ,
    \new_Sorter100|14360_ , \new_Sorter100|14361_ , \new_Sorter100|14362_ ,
    \new_Sorter100|14363_ , \new_Sorter100|14364_ , \new_Sorter100|14365_ ,
    \new_Sorter100|14366_ , \new_Sorter100|14367_ , \new_Sorter100|14368_ ,
    \new_Sorter100|14369_ , \new_Sorter100|14370_ , \new_Sorter100|14371_ ,
    \new_Sorter100|14372_ , \new_Sorter100|14373_ , \new_Sorter100|14374_ ,
    \new_Sorter100|14375_ , \new_Sorter100|14376_ , \new_Sorter100|14377_ ,
    \new_Sorter100|14378_ , \new_Sorter100|14379_ , \new_Sorter100|14380_ ,
    \new_Sorter100|14381_ , \new_Sorter100|14382_ , \new_Sorter100|14383_ ,
    \new_Sorter100|14384_ , \new_Sorter100|14385_ , \new_Sorter100|14386_ ,
    \new_Sorter100|14387_ , \new_Sorter100|14388_ , \new_Sorter100|14389_ ,
    \new_Sorter100|14390_ , \new_Sorter100|14391_ , \new_Sorter100|14392_ ,
    \new_Sorter100|14393_ , \new_Sorter100|14394_ , \new_Sorter100|14395_ ,
    \new_Sorter100|14396_ , \new_Sorter100|14397_ , \new_Sorter100|14398_ ,
    \new_Sorter100|14400_ , \new_Sorter100|14401_ , \new_Sorter100|14402_ ,
    \new_Sorter100|14403_ , \new_Sorter100|14404_ , \new_Sorter100|14405_ ,
    \new_Sorter100|14406_ , \new_Sorter100|14407_ , \new_Sorter100|14408_ ,
    \new_Sorter100|14409_ , \new_Sorter100|14410_ , \new_Sorter100|14411_ ,
    \new_Sorter100|14412_ , \new_Sorter100|14413_ , \new_Sorter100|14414_ ,
    \new_Sorter100|14415_ , \new_Sorter100|14416_ , \new_Sorter100|14417_ ,
    \new_Sorter100|14418_ , \new_Sorter100|14419_ , \new_Sorter100|14420_ ,
    \new_Sorter100|14421_ , \new_Sorter100|14422_ , \new_Sorter100|14423_ ,
    \new_Sorter100|14424_ , \new_Sorter100|14425_ , \new_Sorter100|14426_ ,
    \new_Sorter100|14427_ , \new_Sorter100|14428_ , \new_Sorter100|14429_ ,
    \new_Sorter100|14430_ , \new_Sorter100|14431_ , \new_Sorter100|14432_ ,
    \new_Sorter100|14433_ , \new_Sorter100|14434_ , \new_Sorter100|14435_ ,
    \new_Sorter100|14436_ , \new_Sorter100|14437_ , \new_Sorter100|14438_ ,
    \new_Sorter100|14439_ , \new_Sorter100|14440_ , \new_Sorter100|14441_ ,
    \new_Sorter100|14442_ , \new_Sorter100|14443_ , \new_Sorter100|14444_ ,
    \new_Sorter100|14445_ , \new_Sorter100|14446_ , \new_Sorter100|14447_ ,
    \new_Sorter100|14448_ , \new_Sorter100|14449_ , \new_Sorter100|14450_ ,
    \new_Sorter100|14451_ , \new_Sorter100|14452_ , \new_Sorter100|14453_ ,
    \new_Sorter100|14454_ , \new_Sorter100|14455_ , \new_Sorter100|14456_ ,
    \new_Sorter100|14457_ , \new_Sorter100|14458_ , \new_Sorter100|14459_ ,
    \new_Sorter100|14460_ , \new_Sorter100|14461_ , \new_Sorter100|14462_ ,
    \new_Sorter100|14463_ , \new_Sorter100|14464_ , \new_Sorter100|14465_ ,
    \new_Sorter100|14466_ , \new_Sorter100|14467_ , \new_Sorter100|14468_ ,
    \new_Sorter100|14469_ , \new_Sorter100|14470_ , \new_Sorter100|14471_ ,
    \new_Sorter100|14472_ , \new_Sorter100|14473_ , \new_Sorter100|14474_ ,
    \new_Sorter100|14475_ , \new_Sorter100|14476_ , \new_Sorter100|14477_ ,
    \new_Sorter100|14478_ , \new_Sorter100|14479_ , \new_Sorter100|14480_ ,
    \new_Sorter100|14481_ , \new_Sorter100|14482_ , \new_Sorter100|14483_ ,
    \new_Sorter100|14484_ , \new_Sorter100|14485_ , \new_Sorter100|14486_ ,
    \new_Sorter100|14487_ , \new_Sorter100|14488_ , \new_Sorter100|14489_ ,
    \new_Sorter100|14490_ , \new_Sorter100|14491_ , \new_Sorter100|14492_ ,
    \new_Sorter100|14493_ , \new_Sorter100|14494_ , \new_Sorter100|14495_ ,
    \new_Sorter100|14496_ , \new_Sorter100|14497_ , \new_Sorter100|14498_ ,
    \new_Sorter100|14499_ , \new_Sorter100|14500_ , \new_Sorter100|14599_ ,
    \new_Sorter100|14501_ , \new_Sorter100|14502_ , \new_Sorter100|14503_ ,
    \new_Sorter100|14504_ , \new_Sorter100|14505_ , \new_Sorter100|14506_ ,
    \new_Sorter100|14507_ , \new_Sorter100|14508_ , \new_Sorter100|14509_ ,
    \new_Sorter100|14510_ , \new_Sorter100|14511_ , \new_Sorter100|14512_ ,
    \new_Sorter100|14513_ , \new_Sorter100|14514_ , \new_Sorter100|14515_ ,
    \new_Sorter100|14516_ , \new_Sorter100|14517_ , \new_Sorter100|14518_ ,
    \new_Sorter100|14519_ , \new_Sorter100|14520_ , \new_Sorter100|14521_ ,
    \new_Sorter100|14522_ , \new_Sorter100|14523_ , \new_Sorter100|14524_ ,
    \new_Sorter100|14525_ , \new_Sorter100|14526_ , \new_Sorter100|14527_ ,
    \new_Sorter100|14528_ , \new_Sorter100|14529_ , \new_Sorter100|14530_ ,
    \new_Sorter100|14531_ , \new_Sorter100|14532_ , \new_Sorter100|14533_ ,
    \new_Sorter100|14534_ , \new_Sorter100|14535_ , \new_Sorter100|14536_ ,
    \new_Sorter100|14537_ , \new_Sorter100|14538_ , \new_Sorter100|14539_ ,
    \new_Sorter100|14540_ , \new_Sorter100|14541_ , \new_Sorter100|14542_ ,
    \new_Sorter100|14543_ , \new_Sorter100|14544_ , \new_Sorter100|14545_ ,
    \new_Sorter100|14546_ , \new_Sorter100|14547_ , \new_Sorter100|14548_ ,
    \new_Sorter100|14549_ , \new_Sorter100|14550_ , \new_Sorter100|14551_ ,
    \new_Sorter100|14552_ , \new_Sorter100|14553_ , \new_Sorter100|14554_ ,
    \new_Sorter100|14555_ , \new_Sorter100|14556_ , \new_Sorter100|14557_ ,
    \new_Sorter100|14558_ , \new_Sorter100|14559_ , \new_Sorter100|14560_ ,
    \new_Sorter100|14561_ , \new_Sorter100|14562_ , \new_Sorter100|14563_ ,
    \new_Sorter100|14564_ , \new_Sorter100|14565_ , \new_Sorter100|14566_ ,
    \new_Sorter100|14567_ , \new_Sorter100|14568_ , \new_Sorter100|14569_ ,
    \new_Sorter100|14570_ , \new_Sorter100|14571_ , \new_Sorter100|14572_ ,
    \new_Sorter100|14573_ , \new_Sorter100|14574_ , \new_Sorter100|14575_ ,
    \new_Sorter100|14576_ , \new_Sorter100|14577_ , \new_Sorter100|14578_ ,
    \new_Sorter100|14579_ , \new_Sorter100|14580_ , \new_Sorter100|14581_ ,
    \new_Sorter100|14582_ , \new_Sorter100|14583_ , \new_Sorter100|14584_ ,
    \new_Sorter100|14585_ , \new_Sorter100|14586_ , \new_Sorter100|14587_ ,
    \new_Sorter100|14588_ , \new_Sorter100|14589_ , \new_Sorter100|14590_ ,
    \new_Sorter100|14591_ , \new_Sorter100|14592_ , \new_Sorter100|14593_ ,
    \new_Sorter100|14594_ , \new_Sorter100|14595_ , \new_Sorter100|14596_ ,
    \new_Sorter100|14597_ , \new_Sorter100|14598_ , \new_Sorter100|14600_ ,
    \new_Sorter100|14601_ , \new_Sorter100|14602_ , \new_Sorter100|14603_ ,
    \new_Sorter100|14604_ , \new_Sorter100|14605_ , \new_Sorter100|14606_ ,
    \new_Sorter100|14607_ , \new_Sorter100|14608_ , \new_Sorter100|14609_ ,
    \new_Sorter100|14610_ , \new_Sorter100|14611_ , \new_Sorter100|14612_ ,
    \new_Sorter100|14613_ , \new_Sorter100|14614_ , \new_Sorter100|14615_ ,
    \new_Sorter100|14616_ , \new_Sorter100|14617_ , \new_Sorter100|14618_ ,
    \new_Sorter100|14619_ , \new_Sorter100|14620_ , \new_Sorter100|14621_ ,
    \new_Sorter100|14622_ , \new_Sorter100|14623_ , \new_Sorter100|14624_ ,
    \new_Sorter100|14625_ , \new_Sorter100|14626_ , \new_Sorter100|14627_ ,
    \new_Sorter100|14628_ , \new_Sorter100|14629_ , \new_Sorter100|14630_ ,
    \new_Sorter100|14631_ , \new_Sorter100|14632_ , \new_Sorter100|14633_ ,
    \new_Sorter100|14634_ , \new_Sorter100|14635_ , \new_Sorter100|14636_ ,
    \new_Sorter100|14637_ , \new_Sorter100|14638_ , \new_Sorter100|14639_ ,
    \new_Sorter100|14640_ , \new_Sorter100|14641_ , \new_Sorter100|14642_ ,
    \new_Sorter100|14643_ , \new_Sorter100|14644_ , \new_Sorter100|14645_ ,
    \new_Sorter100|14646_ , \new_Sorter100|14647_ , \new_Sorter100|14648_ ,
    \new_Sorter100|14649_ , \new_Sorter100|14650_ , \new_Sorter100|14651_ ,
    \new_Sorter100|14652_ , \new_Sorter100|14653_ , \new_Sorter100|14654_ ,
    \new_Sorter100|14655_ , \new_Sorter100|14656_ , \new_Sorter100|14657_ ,
    \new_Sorter100|14658_ , \new_Sorter100|14659_ , \new_Sorter100|14660_ ,
    \new_Sorter100|14661_ , \new_Sorter100|14662_ , \new_Sorter100|14663_ ,
    \new_Sorter100|14664_ , \new_Sorter100|14665_ , \new_Sorter100|14666_ ,
    \new_Sorter100|14667_ , \new_Sorter100|14668_ , \new_Sorter100|14669_ ,
    \new_Sorter100|14670_ , \new_Sorter100|14671_ , \new_Sorter100|14672_ ,
    \new_Sorter100|14673_ , \new_Sorter100|14674_ , \new_Sorter100|14675_ ,
    \new_Sorter100|14676_ , \new_Sorter100|14677_ , \new_Sorter100|14678_ ,
    \new_Sorter100|14679_ , \new_Sorter100|14680_ , \new_Sorter100|14681_ ,
    \new_Sorter100|14682_ , \new_Sorter100|14683_ , \new_Sorter100|14684_ ,
    \new_Sorter100|14685_ , \new_Sorter100|14686_ , \new_Sorter100|14687_ ,
    \new_Sorter100|14688_ , \new_Sorter100|14689_ , \new_Sorter100|14690_ ,
    \new_Sorter100|14691_ , \new_Sorter100|14692_ , \new_Sorter100|14693_ ,
    \new_Sorter100|14694_ , \new_Sorter100|14695_ , \new_Sorter100|14696_ ,
    \new_Sorter100|14697_ , \new_Sorter100|14698_ , \new_Sorter100|14699_ ,
    \new_Sorter100|14700_ , \new_Sorter100|14799_ , \new_Sorter100|14701_ ,
    \new_Sorter100|14702_ , \new_Sorter100|14703_ , \new_Sorter100|14704_ ,
    \new_Sorter100|14705_ , \new_Sorter100|14706_ , \new_Sorter100|14707_ ,
    \new_Sorter100|14708_ , \new_Sorter100|14709_ , \new_Sorter100|14710_ ,
    \new_Sorter100|14711_ , \new_Sorter100|14712_ , \new_Sorter100|14713_ ,
    \new_Sorter100|14714_ , \new_Sorter100|14715_ , \new_Sorter100|14716_ ,
    \new_Sorter100|14717_ , \new_Sorter100|14718_ , \new_Sorter100|14719_ ,
    \new_Sorter100|14720_ , \new_Sorter100|14721_ , \new_Sorter100|14722_ ,
    \new_Sorter100|14723_ , \new_Sorter100|14724_ , \new_Sorter100|14725_ ,
    \new_Sorter100|14726_ , \new_Sorter100|14727_ , \new_Sorter100|14728_ ,
    \new_Sorter100|14729_ , \new_Sorter100|14730_ , \new_Sorter100|14731_ ,
    \new_Sorter100|14732_ , \new_Sorter100|14733_ , \new_Sorter100|14734_ ,
    \new_Sorter100|14735_ , \new_Sorter100|14736_ , \new_Sorter100|14737_ ,
    \new_Sorter100|14738_ , \new_Sorter100|14739_ , \new_Sorter100|14740_ ,
    \new_Sorter100|14741_ , \new_Sorter100|14742_ , \new_Sorter100|14743_ ,
    \new_Sorter100|14744_ , \new_Sorter100|14745_ , \new_Sorter100|14746_ ,
    \new_Sorter100|14747_ , \new_Sorter100|14748_ , \new_Sorter100|14749_ ,
    \new_Sorter100|14750_ , \new_Sorter100|14751_ , \new_Sorter100|14752_ ,
    \new_Sorter100|14753_ , \new_Sorter100|14754_ , \new_Sorter100|14755_ ,
    \new_Sorter100|14756_ , \new_Sorter100|14757_ , \new_Sorter100|14758_ ,
    \new_Sorter100|14759_ , \new_Sorter100|14760_ , \new_Sorter100|14761_ ,
    \new_Sorter100|14762_ , \new_Sorter100|14763_ , \new_Sorter100|14764_ ,
    \new_Sorter100|14765_ , \new_Sorter100|14766_ , \new_Sorter100|14767_ ,
    \new_Sorter100|14768_ , \new_Sorter100|14769_ , \new_Sorter100|14770_ ,
    \new_Sorter100|14771_ , \new_Sorter100|14772_ , \new_Sorter100|14773_ ,
    \new_Sorter100|14774_ , \new_Sorter100|14775_ , \new_Sorter100|14776_ ,
    \new_Sorter100|14777_ , \new_Sorter100|14778_ , \new_Sorter100|14779_ ,
    \new_Sorter100|14780_ , \new_Sorter100|14781_ , \new_Sorter100|14782_ ,
    \new_Sorter100|14783_ , \new_Sorter100|14784_ , \new_Sorter100|14785_ ,
    \new_Sorter100|14786_ , \new_Sorter100|14787_ , \new_Sorter100|14788_ ,
    \new_Sorter100|14789_ , \new_Sorter100|14790_ , \new_Sorter100|14791_ ,
    \new_Sorter100|14792_ , \new_Sorter100|14793_ , \new_Sorter100|14794_ ,
    \new_Sorter100|14795_ , \new_Sorter100|14796_ , \new_Sorter100|14797_ ,
    \new_Sorter100|14798_ , \new_Sorter100|14800_ , \new_Sorter100|14801_ ,
    \new_Sorter100|14802_ , \new_Sorter100|14803_ , \new_Sorter100|14804_ ,
    \new_Sorter100|14805_ , \new_Sorter100|14806_ , \new_Sorter100|14807_ ,
    \new_Sorter100|14808_ , \new_Sorter100|14809_ , \new_Sorter100|14810_ ,
    \new_Sorter100|14811_ , \new_Sorter100|14812_ , \new_Sorter100|14813_ ,
    \new_Sorter100|14814_ , \new_Sorter100|14815_ , \new_Sorter100|14816_ ,
    \new_Sorter100|14817_ , \new_Sorter100|14818_ , \new_Sorter100|14819_ ,
    \new_Sorter100|14820_ , \new_Sorter100|14821_ , \new_Sorter100|14822_ ,
    \new_Sorter100|14823_ , \new_Sorter100|14824_ , \new_Sorter100|14825_ ,
    \new_Sorter100|14826_ , \new_Sorter100|14827_ , \new_Sorter100|14828_ ,
    \new_Sorter100|14829_ , \new_Sorter100|14830_ , \new_Sorter100|14831_ ,
    \new_Sorter100|14832_ , \new_Sorter100|14833_ , \new_Sorter100|14834_ ,
    \new_Sorter100|14835_ , \new_Sorter100|14836_ , \new_Sorter100|14837_ ,
    \new_Sorter100|14838_ , \new_Sorter100|14839_ , \new_Sorter100|14840_ ,
    \new_Sorter100|14841_ , \new_Sorter100|14842_ , \new_Sorter100|14843_ ,
    \new_Sorter100|14844_ , \new_Sorter100|14845_ , \new_Sorter100|14846_ ,
    \new_Sorter100|14847_ , \new_Sorter100|14848_ , \new_Sorter100|14849_ ,
    \new_Sorter100|14850_ , \new_Sorter100|14851_ , \new_Sorter100|14852_ ,
    \new_Sorter100|14853_ , \new_Sorter100|14854_ , \new_Sorter100|14855_ ,
    \new_Sorter100|14856_ , \new_Sorter100|14857_ , \new_Sorter100|14858_ ,
    \new_Sorter100|14859_ , \new_Sorter100|14860_ , \new_Sorter100|14861_ ,
    \new_Sorter100|14862_ , \new_Sorter100|14863_ , \new_Sorter100|14864_ ,
    \new_Sorter100|14865_ , \new_Sorter100|14866_ , \new_Sorter100|14867_ ,
    \new_Sorter100|14868_ , \new_Sorter100|14869_ , \new_Sorter100|14870_ ,
    \new_Sorter100|14871_ , \new_Sorter100|14872_ , \new_Sorter100|14873_ ,
    \new_Sorter100|14874_ , \new_Sorter100|14875_ , \new_Sorter100|14876_ ,
    \new_Sorter100|14877_ , \new_Sorter100|14878_ , \new_Sorter100|14879_ ,
    \new_Sorter100|14880_ , \new_Sorter100|14881_ , \new_Sorter100|14882_ ,
    \new_Sorter100|14883_ , \new_Sorter100|14884_ , \new_Sorter100|14885_ ,
    \new_Sorter100|14886_ , \new_Sorter100|14887_ , \new_Sorter100|14888_ ,
    \new_Sorter100|14889_ , \new_Sorter100|14890_ , \new_Sorter100|14891_ ,
    \new_Sorter100|14892_ , \new_Sorter100|14893_ , \new_Sorter100|14894_ ,
    \new_Sorter100|14895_ , \new_Sorter100|14896_ , \new_Sorter100|14897_ ,
    \new_Sorter100|14898_ , \new_Sorter100|14899_ , \new_Sorter100|14900_ ,
    \new_Sorter100|14999_ , \new_Sorter100|14901_ , \new_Sorter100|14902_ ,
    \new_Sorter100|14903_ , \new_Sorter100|14904_ , \new_Sorter100|14905_ ,
    \new_Sorter100|14906_ , \new_Sorter100|14907_ , \new_Sorter100|14908_ ,
    \new_Sorter100|14909_ , \new_Sorter100|14910_ , \new_Sorter100|14911_ ,
    \new_Sorter100|14912_ , \new_Sorter100|14913_ , \new_Sorter100|14914_ ,
    \new_Sorter100|14915_ , \new_Sorter100|14916_ , \new_Sorter100|14917_ ,
    \new_Sorter100|14918_ , \new_Sorter100|14919_ , \new_Sorter100|14920_ ,
    \new_Sorter100|14921_ , \new_Sorter100|14922_ , \new_Sorter100|14923_ ,
    \new_Sorter100|14924_ , \new_Sorter100|14925_ , \new_Sorter100|14926_ ,
    \new_Sorter100|14927_ , \new_Sorter100|14928_ , \new_Sorter100|14929_ ,
    \new_Sorter100|14930_ , \new_Sorter100|14931_ , \new_Sorter100|14932_ ,
    \new_Sorter100|14933_ , \new_Sorter100|14934_ , \new_Sorter100|14935_ ,
    \new_Sorter100|14936_ , \new_Sorter100|14937_ , \new_Sorter100|14938_ ,
    \new_Sorter100|14939_ , \new_Sorter100|14940_ , \new_Sorter100|14941_ ,
    \new_Sorter100|14942_ , \new_Sorter100|14943_ , \new_Sorter100|14944_ ,
    \new_Sorter100|14945_ , \new_Sorter100|14946_ , \new_Sorter100|14947_ ,
    \new_Sorter100|14948_ , \new_Sorter100|14949_ , \new_Sorter100|14950_ ,
    \new_Sorter100|14951_ , \new_Sorter100|14952_ , \new_Sorter100|14953_ ,
    \new_Sorter100|14954_ , \new_Sorter100|14955_ , \new_Sorter100|14956_ ,
    \new_Sorter100|14957_ , \new_Sorter100|14958_ , \new_Sorter100|14959_ ,
    \new_Sorter100|14960_ , \new_Sorter100|14961_ , \new_Sorter100|14962_ ,
    \new_Sorter100|14963_ , \new_Sorter100|14964_ , \new_Sorter100|14965_ ,
    \new_Sorter100|14966_ , \new_Sorter100|14967_ , \new_Sorter100|14968_ ,
    \new_Sorter100|14969_ , \new_Sorter100|14970_ , \new_Sorter100|14971_ ,
    \new_Sorter100|14972_ , \new_Sorter100|14973_ , \new_Sorter100|14974_ ,
    \new_Sorter100|14975_ , \new_Sorter100|14976_ , \new_Sorter100|14977_ ,
    \new_Sorter100|14978_ , \new_Sorter100|14979_ , \new_Sorter100|14980_ ,
    \new_Sorter100|14981_ , \new_Sorter100|14982_ , \new_Sorter100|14983_ ,
    \new_Sorter100|14984_ , \new_Sorter100|14985_ , \new_Sorter100|14986_ ,
    \new_Sorter100|14987_ , \new_Sorter100|14988_ , \new_Sorter100|14989_ ,
    \new_Sorter100|14990_ , \new_Sorter100|14991_ , \new_Sorter100|14992_ ,
    \new_Sorter100|14993_ , \new_Sorter100|14994_ , \new_Sorter100|14995_ ,
    \new_Sorter100|14996_ , \new_Sorter100|14997_ , \new_Sorter100|14998_ ,
    \new_Sorter100|15000_ , \new_Sorter100|15001_ , \new_Sorter100|15002_ ,
    \new_Sorter100|15003_ , \new_Sorter100|15004_ , \new_Sorter100|15005_ ,
    \new_Sorter100|15006_ , \new_Sorter100|15007_ , \new_Sorter100|15008_ ,
    \new_Sorter100|15009_ , \new_Sorter100|15010_ , \new_Sorter100|15011_ ,
    \new_Sorter100|15012_ , \new_Sorter100|15013_ , \new_Sorter100|15014_ ,
    \new_Sorter100|15015_ , \new_Sorter100|15016_ , \new_Sorter100|15017_ ,
    \new_Sorter100|15018_ , \new_Sorter100|15019_ , \new_Sorter100|15020_ ,
    \new_Sorter100|15021_ , \new_Sorter100|15022_ , \new_Sorter100|15023_ ,
    \new_Sorter100|15024_ , \new_Sorter100|15025_ , \new_Sorter100|15026_ ,
    \new_Sorter100|15027_ , \new_Sorter100|15028_ , \new_Sorter100|15029_ ,
    \new_Sorter100|15030_ , \new_Sorter100|15031_ , \new_Sorter100|15032_ ,
    \new_Sorter100|15033_ , \new_Sorter100|15034_ , \new_Sorter100|15035_ ,
    \new_Sorter100|15036_ , \new_Sorter100|15037_ , \new_Sorter100|15038_ ,
    \new_Sorter100|15039_ , \new_Sorter100|15040_ , \new_Sorter100|15041_ ,
    \new_Sorter100|15042_ , \new_Sorter100|15043_ , \new_Sorter100|15044_ ,
    \new_Sorter100|15045_ , \new_Sorter100|15046_ , \new_Sorter100|15047_ ,
    \new_Sorter100|15048_ , \new_Sorter100|15049_ , \new_Sorter100|15050_ ,
    \new_Sorter100|15051_ , \new_Sorter100|15052_ , \new_Sorter100|15053_ ,
    \new_Sorter100|15054_ , \new_Sorter100|15055_ , \new_Sorter100|15056_ ,
    \new_Sorter100|15057_ , \new_Sorter100|15058_ , \new_Sorter100|15059_ ,
    \new_Sorter100|15060_ , \new_Sorter100|15061_ , \new_Sorter100|15062_ ,
    \new_Sorter100|15063_ , \new_Sorter100|15064_ , \new_Sorter100|15065_ ,
    \new_Sorter100|15066_ , \new_Sorter100|15067_ , \new_Sorter100|15068_ ,
    \new_Sorter100|15069_ , \new_Sorter100|15070_ , \new_Sorter100|15071_ ,
    \new_Sorter100|15072_ , \new_Sorter100|15073_ , \new_Sorter100|15074_ ,
    \new_Sorter100|15075_ , \new_Sorter100|15076_ , \new_Sorter100|15077_ ,
    \new_Sorter100|15078_ , \new_Sorter100|15079_ , \new_Sorter100|15080_ ,
    \new_Sorter100|15081_ , \new_Sorter100|15082_ , \new_Sorter100|15083_ ,
    \new_Sorter100|15084_ , \new_Sorter100|15085_ , \new_Sorter100|15086_ ,
    \new_Sorter100|15087_ , \new_Sorter100|15088_ , \new_Sorter100|15089_ ,
    \new_Sorter100|15090_ , \new_Sorter100|15091_ , \new_Sorter100|15092_ ,
    \new_Sorter100|15093_ , \new_Sorter100|15094_ , \new_Sorter100|15095_ ,
    \new_Sorter100|15096_ , \new_Sorter100|15097_ , \new_Sorter100|15098_ ,
    \new_Sorter100|15099_ , \new_Sorter100|15100_ , \new_Sorter100|15199_ ,
    \new_Sorter100|15101_ , \new_Sorter100|15102_ , \new_Sorter100|15103_ ,
    \new_Sorter100|15104_ , \new_Sorter100|15105_ , \new_Sorter100|15106_ ,
    \new_Sorter100|15107_ , \new_Sorter100|15108_ , \new_Sorter100|15109_ ,
    \new_Sorter100|15110_ , \new_Sorter100|15111_ , \new_Sorter100|15112_ ,
    \new_Sorter100|15113_ , \new_Sorter100|15114_ , \new_Sorter100|15115_ ,
    \new_Sorter100|15116_ , \new_Sorter100|15117_ , \new_Sorter100|15118_ ,
    \new_Sorter100|15119_ , \new_Sorter100|15120_ , \new_Sorter100|15121_ ,
    \new_Sorter100|15122_ , \new_Sorter100|15123_ , \new_Sorter100|15124_ ,
    \new_Sorter100|15125_ , \new_Sorter100|15126_ , \new_Sorter100|15127_ ,
    \new_Sorter100|15128_ , \new_Sorter100|15129_ , \new_Sorter100|15130_ ,
    \new_Sorter100|15131_ , \new_Sorter100|15132_ , \new_Sorter100|15133_ ,
    \new_Sorter100|15134_ , \new_Sorter100|15135_ , \new_Sorter100|15136_ ,
    \new_Sorter100|15137_ , \new_Sorter100|15138_ , \new_Sorter100|15139_ ,
    \new_Sorter100|15140_ , \new_Sorter100|15141_ , \new_Sorter100|15142_ ,
    \new_Sorter100|15143_ , \new_Sorter100|15144_ , \new_Sorter100|15145_ ,
    \new_Sorter100|15146_ , \new_Sorter100|15147_ , \new_Sorter100|15148_ ,
    \new_Sorter100|15149_ , \new_Sorter100|15150_ , \new_Sorter100|15151_ ,
    \new_Sorter100|15152_ , \new_Sorter100|15153_ , \new_Sorter100|15154_ ,
    \new_Sorter100|15155_ , \new_Sorter100|15156_ , \new_Sorter100|15157_ ,
    \new_Sorter100|15158_ , \new_Sorter100|15159_ , \new_Sorter100|15160_ ,
    \new_Sorter100|15161_ , \new_Sorter100|15162_ , \new_Sorter100|15163_ ,
    \new_Sorter100|15164_ , \new_Sorter100|15165_ , \new_Sorter100|15166_ ,
    \new_Sorter100|15167_ , \new_Sorter100|15168_ , \new_Sorter100|15169_ ,
    \new_Sorter100|15170_ , \new_Sorter100|15171_ , \new_Sorter100|15172_ ,
    \new_Sorter100|15173_ , \new_Sorter100|15174_ , \new_Sorter100|15175_ ,
    \new_Sorter100|15176_ , \new_Sorter100|15177_ , \new_Sorter100|15178_ ,
    \new_Sorter100|15179_ , \new_Sorter100|15180_ , \new_Sorter100|15181_ ,
    \new_Sorter100|15182_ , \new_Sorter100|15183_ , \new_Sorter100|15184_ ,
    \new_Sorter100|15185_ , \new_Sorter100|15186_ , \new_Sorter100|15187_ ,
    \new_Sorter100|15188_ , \new_Sorter100|15189_ , \new_Sorter100|15190_ ,
    \new_Sorter100|15191_ , \new_Sorter100|15192_ , \new_Sorter100|15193_ ,
    \new_Sorter100|15194_ , \new_Sorter100|15195_ , \new_Sorter100|15196_ ,
    \new_Sorter100|15197_ , \new_Sorter100|15198_ , \new_Sorter100|15200_ ,
    \new_Sorter100|15201_ , \new_Sorter100|15202_ , \new_Sorter100|15203_ ,
    \new_Sorter100|15204_ , \new_Sorter100|15205_ , \new_Sorter100|15206_ ,
    \new_Sorter100|15207_ , \new_Sorter100|15208_ , \new_Sorter100|15209_ ,
    \new_Sorter100|15210_ , \new_Sorter100|15211_ , \new_Sorter100|15212_ ,
    \new_Sorter100|15213_ , \new_Sorter100|15214_ , \new_Sorter100|15215_ ,
    \new_Sorter100|15216_ , \new_Sorter100|15217_ , \new_Sorter100|15218_ ,
    \new_Sorter100|15219_ , \new_Sorter100|15220_ , \new_Sorter100|15221_ ,
    \new_Sorter100|15222_ , \new_Sorter100|15223_ , \new_Sorter100|15224_ ,
    \new_Sorter100|15225_ , \new_Sorter100|15226_ , \new_Sorter100|15227_ ,
    \new_Sorter100|15228_ , \new_Sorter100|15229_ , \new_Sorter100|15230_ ,
    \new_Sorter100|15231_ , \new_Sorter100|15232_ , \new_Sorter100|15233_ ,
    \new_Sorter100|15234_ , \new_Sorter100|15235_ , \new_Sorter100|15236_ ,
    \new_Sorter100|15237_ , \new_Sorter100|15238_ , \new_Sorter100|15239_ ,
    \new_Sorter100|15240_ , \new_Sorter100|15241_ , \new_Sorter100|15242_ ,
    \new_Sorter100|15243_ , \new_Sorter100|15244_ , \new_Sorter100|15245_ ,
    \new_Sorter100|15246_ , \new_Sorter100|15247_ , \new_Sorter100|15248_ ,
    \new_Sorter100|15249_ , \new_Sorter100|15250_ , \new_Sorter100|15251_ ,
    \new_Sorter100|15252_ , \new_Sorter100|15253_ , \new_Sorter100|15254_ ,
    \new_Sorter100|15255_ , \new_Sorter100|15256_ , \new_Sorter100|15257_ ,
    \new_Sorter100|15258_ , \new_Sorter100|15259_ , \new_Sorter100|15260_ ,
    \new_Sorter100|15261_ , \new_Sorter100|15262_ , \new_Sorter100|15263_ ,
    \new_Sorter100|15264_ , \new_Sorter100|15265_ , \new_Sorter100|15266_ ,
    \new_Sorter100|15267_ , \new_Sorter100|15268_ , \new_Sorter100|15269_ ,
    \new_Sorter100|15270_ , \new_Sorter100|15271_ , \new_Sorter100|15272_ ,
    \new_Sorter100|15273_ , \new_Sorter100|15274_ , \new_Sorter100|15275_ ,
    \new_Sorter100|15276_ , \new_Sorter100|15277_ , \new_Sorter100|15278_ ,
    \new_Sorter100|15279_ , \new_Sorter100|15280_ , \new_Sorter100|15281_ ,
    \new_Sorter100|15282_ , \new_Sorter100|15283_ , \new_Sorter100|15284_ ,
    \new_Sorter100|15285_ , \new_Sorter100|15286_ , \new_Sorter100|15287_ ,
    \new_Sorter100|15288_ , \new_Sorter100|15289_ , \new_Sorter100|15290_ ,
    \new_Sorter100|15291_ , \new_Sorter100|15292_ , \new_Sorter100|15293_ ,
    \new_Sorter100|15294_ , \new_Sorter100|15295_ , \new_Sorter100|15296_ ,
    \new_Sorter100|15297_ , \new_Sorter100|15298_ , \new_Sorter100|15299_ ,
    \new_Sorter100|15300_ , \new_Sorter100|15399_ , \new_Sorter100|15301_ ,
    \new_Sorter100|15302_ , \new_Sorter100|15303_ , \new_Sorter100|15304_ ,
    \new_Sorter100|15305_ , \new_Sorter100|15306_ , \new_Sorter100|15307_ ,
    \new_Sorter100|15308_ , \new_Sorter100|15309_ , \new_Sorter100|15310_ ,
    \new_Sorter100|15311_ , \new_Sorter100|15312_ , \new_Sorter100|15313_ ,
    \new_Sorter100|15314_ , \new_Sorter100|15315_ , \new_Sorter100|15316_ ,
    \new_Sorter100|15317_ , \new_Sorter100|15318_ , \new_Sorter100|15319_ ,
    \new_Sorter100|15320_ , \new_Sorter100|15321_ , \new_Sorter100|15322_ ,
    \new_Sorter100|15323_ , \new_Sorter100|15324_ , \new_Sorter100|15325_ ,
    \new_Sorter100|15326_ , \new_Sorter100|15327_ , \new_Sorter100|15328_ ,
    \new_Sorter100|15329_ , \new_Sorter100|15330_ , \new_Sorter100|15331_ ,
    \new_Sorter100|15332_ , \new_Sorter100|15333_ , \new_Sorter100|15334_ ,
    \new_Sorter100|15335_ , \new_Sorter100|15336_ , \new_Sorter100|15337_ ,
    \new_Sorter100|15338_ , \new_Sorter100|15339_ , \new_Sorter100|15340_ ,
    \new_Sorter100|15341_ , \new_Sorter100|15342_ , \new_Sorter100|15343_ ,
    \new_Sorter100|15344_ , \new_Sorter100|15345_ , \new_Sorter100|15346_ ,
    \new_Sorter100|15347_ , \new_Sorter100|15348_ , \new_Sorter100|15349_ ,
    \new_Sorter100|15350_ , \new_Sorter100|15351_ , \new_Sorter100|15352_ ,
    \new_Sorter100|15353_ , \new_Sorter100|15354_ , \new_Sorter100|15355_ ,
    \new_Sorter100|15356_ , \new_Sorter100|15357_ , \new_Sorter100|15358_ ,
    \new_Sorter100|15359_ , \new_Sorter100|15360_ , \new_Sorter100|15361_ ,
    \new_Sorter100|15362_ , \new_Sorter100|15363_ , \new_Sorter100|15364_ ,
    \new_Sorter100|15365_ , \new_Sorter100|15366_ , \new_Sorter100|15367_ ,
    \new_Sorter100|15368_ , \new_Sorter100|15369_ , \new_Sorter100|15370_ ,
    \new_Sorter100|15371_ , \new_Sorter100|15372_ , \new_Sorter100|15373_ ,
    \new_Sorter100|15374_ , \new_Sorter100|15375_ , \new_Sorter100|15376_ ,
    \new_Sorter100|15377_ , \new_Sorter100|15378_ , \new_Sorter100|15379_ ,
    \new_Sorter100|15380_ , \new_Sorter100|15381_ , \new_Sorter100|15382_ ,
    \new_Sorter100|15383_ , \new_Sorter100|15384_ , \new_Sorter100|15385_ ,
    \new_Sorter100|15386_ , \new_Sorter100|15387_ , \new_Sorter100|15388_ ,
    \new_Sorter100|15389_ , \new_Sorter100|15390_ , \new_Sorter100|15391_ ,
    \new_Sorter100|15392_ , \new_Sorter100|15393_ , \new_Sorter100|15394_ ,
    \new_Sorter100|15395_ , \new_Sorter100|15396_ , \new_Sorter100|15397_ ,
    \new_Sorter100|15398_ , \new_Sorter100|15400_ , \new_Sorter100|15401_ ,
    \new_Sorter100|15402_ , \new_Sorter100|15403_ , \new_Sorter100|15404_ ,
    \new_Sorter100|15405_ , \new_Sorter100|15406_ , \new_Sorter100|15407_ ,
    \new_Sorter100|15408_ , \new_Sorter100|15409_ , \new_Sorter100|15410_ ,
    \new_Sorter100|15411_ , \new_Sorter100|15412_ , \new_Sorter100|15413_ ,
    \new_Sorter100|15414_ , \new_Sorter100|15415_ , \new_Sorter100|15416_ ,
    \new_Sorter100|15417_ , \new_Sorter100|15418_ , \new_Sorter100|15419_ ,
    \new_Sorter100|15420_ , \new_Sorter100|15421_ , \new_Sorter100|15422_ ,
    \new_Sorter100|15423_ , \new_Sorter100|15424_ , \new_Sorter100|15425_ ,
    \new_Sorter100|15426_ , \new_Sorter100|15427_ , \new_Sorter100|15428_ ,
    \new_Sorter100|15429_ , \new_Sorter100|15430_ , \new_Sorter100|15431_ ,
    \new_Sorter100|15432_ , \new_Sorter100|15433_ , \new_Sorter100|15434_ ,
    \new_Sorter100|15435_ , \new_Sorter100|15436_ , \new_Sorter100|15437_ ,
    \new_Sorter100|15438_ , \new_Sorter100|15439_ , \new_Sorter100|15440_ ,
    \new_Sorter100|15441_ , \new_Sorter100|15442_ , \new_Sorter100|15443_ ,
    \new_Sorter100|15444_ , \new_Sorter100|15445_ , \new_Sorter100|15446_ ,
    \new_Sorter100|15447_ , \new_Sorter100|15448_ , \new_Sorter100|15449_ ,
    \new_Sorter100|15450_ , \new_Sorter100|15451_ , \new_Sorter100|15452_ ,
    \new_Sorter100|15453_ , \new_Sorter100|15454_ , \new_Sorter100|15455_ ,
    \new_Sorter100|15456_ , \new_Sorter100|15457_ , \new_Sorter100|15458_ ,
    \new_Sorter100|15459_ , \new_Sorter100|15460_ , \new_Sorter100|15461_ ,
    \new_Sorter100|15462_ , \new_Sorter100|15463_ , \new_Sorter100|15464_ ,
    \new_Sorter100|15465_ , \new_Sorter100|15466_ , \new_Sorter100|15467_ ,
    \new_Sorter100|15468_ , \new_Sorter100|15469_ , \new_Sorter100|15470_ ,
    \new_Sorter100|15471_ , \new_Sorter100|15472_ , \new_Sorter100|15473_ ,
    \new_Sorter100|15474_ , \new_Sorter100|15475_ , \new_Sorter100|15476_ ,
    \new_Sorter100|15477_ , \new_Sorter100|15478_ , \new_Sorter100|15479_ ,
    \new_Sorter100|15480_ , \new_Sorter100|15481_ , \new_Sorter100|15482_ ,
    \new_Sorter100|15483_ , \new_Sorter100|15484_ , \new_Sorter100|15485_ ,
    \new_Sorter100|15486_ , \new_Sorter100|15487_ , \new_Sorter100|15488_ ,
    \new_Sorter100|15489_ , \new_Sorter100|15490_ , \new_Sorter100|15491_ ,
    \new_Sorter100|15492_ , \new_Sorter100|15493_ , \new_Sorter100|15494_ ,
    \new_Sorter100|15495_ , \new_Sorter100|15496_ , \new_Sorter100|15497_ ,
    \new_Sorter100|15498_ , \new_Sorter100|15499_ , \new_Sorter100|15500_ ,
    \new_Sorter100|15599_ , \new_Sorter100|15501_ , \new_Sorter100|15502_ ,
    \new_Sorter100|15503_ , \new_Sorter100|15504_ , \new_Sorter100|15505_ ,
    \new_Sorter100|15506_ , \new_Sorter100|15507_ , \new_Sorter100|15508_ ,
    \new_Sorter100|15509_ , \new_Sorter100|15510_ , \new_Sorter100|15511_ ,
    \new_Sorter100|15512_ , \new_Sorter100|15513_ , \new_Sorter100|15514_ ,
    \new_Sorter100|15515_ , \new_Sorter100|15516_ , \new_Sorter100|15517_ ,
    \new_Sorter100|15518_ , \new_Sorter100|15519_ , \new_Sorter100|15520_ ,
    \new_Sorter100|15521_ , \new_Sorter100|15522_ , \new_Sorter100|15523_ ,
    \new_Sorter100|15524_ , \new_Sorter100|15525_ , \new_Sorter100|15526_ ,
    \new_Sorter100|15527_ , \new_Sorter100|15528_ , \new_Sorter100|15529_ ,
    \new_Sorter100|15530_ , \new_Sorter100|15531_ , \new_Sorter100|15532_ ,
    \new_Sorter100|15533_ , \new_Sorter100|15534_ , \new_Sorter100|15535_ ,
    \new_Sorter100|15536_ , \new_Sorter100|15537_ , \new_Sorter100|15538_ ,
    \new_Sorter100|15539_ , \new_Sorter100|15540_ , \new_Sorter100|15541_ ,
    \new_Sorter100|15542_ , \new_Sorter100|15543_ , \new_Sorter100|15544_ ,
    \new_Sorter100|15545_ , \new_Sorter100|15546_ , \new_Sorter100|15547_ ,
    \new_Sorter100|15548_ , \new_Sorter100|15549_ , \new_Sorter100|15550_ ,
    \new_Sorter100|15551_ , \new_Sorter100|15552_ , \new_Sorter100|15553_ ,
    \new_Sorter100|15554_ , \new_Sorter100|15555_ , \new_Sorter100|15556_ ,
    \new_Sorter100|15557_ , \new_Sorter100|15558_ , \new_Sorter100|15559_ ,
    \new_Sorter100|15560_ , \new_Sorter100|15561_ , \new_Sorter100|15562_ ,
    \new_Sorter100|15563_ , \new_Sorter100|15564_ , \new_Sorter100|15565_ ,
    \new_Sorter100|15566_ , \new_Sorter100|15567_ , \new_Sorter100|15568_ ,
    \new_Sorter100|15569_ , \new_Sorter100|15570_ , \new_Sorter100|15571_ ,
    \new_Sorter100|15572_ , \new_Sorter100|15573_ , \new_Sorter100|15574_ ,
    \new_Sorter100|15575_ , \new_Sorter100|15576_ , \new_Sorter100|15577_ ,
    \new_Sorter100|15578_ , \new_Sorter100|15579_ , \new_Sorter100|15580_ ,
    \new_Sorter100|15581_ , \new_Sorter100|15582_ , \new_Sorter100|15583_ ,
    \new_Sorter100|15584_ , \new_Sorter100|15585_ , \new_Sorter100|15586_ ,
    \new_Sorter100|15587_ , \new_Sorter100|15588_ , \new_Sorter100|15589_ ,
    \new_Sorter100|15590_ , \new_Sorter100|15591_ , \new_Sorter100|15592_ ,
    \new_Sorter100|15593_ , \new_Sorter100|15594_ , \new_Sorter100|15595_ ,
    \new_Sorter100|15596_ , \new_Sorter100|15597_ , \new_Sorter100|15598_ ,
    \new_Sorter100|15600_ , \new_Sorter100|15601_ , \new_Sorter100|15602_ ,
    \new_Sorter100|15603_ , \new_Sorter100|15604_ , \new_Sorter100|15605_ ,
    \new_Sorter100|15606_ , \new_Sorter100|15607_ , \new_Sorter100|15608_ ,
    \new_Sorter100|15609_ , \new_Sorter100|15610_ , \new_Sorter100|15611_ ,
    \new_Sorter100|15612_ , \new_Sorter100|15613_ , \new_Sorter100|15614_ ,
    \new_Sorter100|15615_ , \new_Sorter100|15616_ , \new_Sorter100|15617_ ,
    \new_Sorter100|15618_ , \new_Sorter100|15619_ , \new_Sorter100|15620_ ,
    \new_Sorter100|15621_ , \new_Sorter100|15622_ , \new_Sorter100|15623_ ,
    \new_Sorter100|15624_ , \new_Sorter100|15625_ , \new_Sorter100|15626_ ,
    \new_Sorter100|15627_ , \new_Sorter100|15628_ , \new_Sorter100|15629_ ,
    \new_Sorter100|15630_ , \new_Sorter100|15631_ , \new_Sorter100|15632_ ,
    \new_Sorter100|15633_ , \new_Sorter100|15634_ , \new_Sorter100|15635_ ,
    \new_Sorter100|15636_ , \new_Sorter100|15637_ , \new_Sorter100|15638_ ,
    \new_Sorter100|15639_ , \new_Sorter100|15640_ , \new_Sorter100|15641_ ,
    \new_Sorter100|15642_ , \new_Sorter100|15643_ , \new_Sorter100|15644_ ,
    \new_Sorter100|15645_ , \new_Sorter100|15646_ , \new_Sorter100|15647_ ,
    \new_Sorter100|15648_ , \new_Sorter100|15649_ , \new_Sorter100|15650_ ,
    \new_Sorter100|15651_ , \new_Sorter100|15652_ , \new_Sorter100|15653_ ,
    \new_Sorter100|15654_ , \new_Sorter100|15655_ , \new_Sorter100|15656_ ,
    \new_Sorter100|15657_ , \new_Sorter100|15658_ , \new_Sorter100|15659_ ,
    \new_Sorter100|15660_ , \new_Sorter100|15661_ , \new_Sorter100|15662_ ,
    \new_Sorter100|15663_ , \new_Sorter100|15664_ , \new_Sorter100|15665_ ,
    \new_Sorter100|15666_ , \new_Sorter100|15667_ , \new_Sorter100|15668_ ,
    \new_Sorter100|15669_ , \new_Sorter100|15670_ , \new_Sorter100|15671_ ,
    \new_Sorter100|15672_ , \new_Sorter100|15673_ , \new_Sorter100|15674_ ,
    \new_Sorter100|15675_ , \new_Sorter100|15676_ , \new_Sorter100|15677_ ,
    \new_Sorter100|15678_ , \new_Sorter100|15679_ , \new_Sorter100|15680_ ,
    \new_Sorter100|15681_ , \new_Sorter100|15682_ , \new_Sorter100|15683_ ,
    \new_Sorter100|15684_ , \new_Sorter100|15685_ , \new_Sorter100|15686_ ,
    \new_Sorter100|15687_ , \new_Sorter100|15688_ , \new_Sorter100|15689_ ,
    \new_Sorter100|15690_ , \new_Sorter100|15691_ , \new_Sorter100|15692_ ,
    \new_Sorter100|15693_ , \new_Sorter100|15694_ , \new_Sorter100|15695_ ,
    \new_Sorter100|15696_ , \new_Sorter100|15697_ , \new_Sorter100|15698_ ,
    \new_Sorter100|15699_ , \new_Sorter100|15700_ , \new_Sorter100|15799_ ,
    \new_Sorter100|15701_ , \new_Sorter100|15702_ , \new_Sorter100|15703_ ,
    \new_Sorter100|15704_ , \new_Sorter100|15705_ , \new_Sorter100|15706_ ,
    \new_Sorter100|15707_ , \new_Sorter100|15708_ , \new_Sorter100|15709_ ,
    \new_Sorter100|15710_ , \new_Sorter100|15711_ , \new_Sorter100|15712_ ,
    \new_Sorter100|15713_ , \new_Sorter100|15714_ , \new_Sorter100|15715_ ,
    \new_Sorter100|15716_ , \new_Sorter100|15717_ , \new_Sorter100|15718_ ,
    \new_Sorter100|15719_ , \new_Sorter100|15720_ , \new_Sorter100|15721_ ,
    \new_Sorter100|15722_ , \new_Sorter100|15723_ , \new_Sorter100|15724_ ,
    \new_Sorter100|15725_ , \new_Sorter100|15726_ , \new_Sorter100|15727_ ,
    \new_Sorter100|15728_ , \new_Sorter100|15729_ , \new_Sorter100|15730_ ,
    \new_Sorter100|15731_ , \new_Sorter100|15732_ , \new_Sorter100|15733_ ,
    \new_Sorter100|15734_ , \new_Sorter100|15735_ , \new_Sorter100|15736_ ,
    \new_Sorter100|15737_ , \new_Sorter100|15738_ , \new_Sorter100|15739_ ,
    \new_Sorter100|15740_ , \new_Sorter100|15741_ , \new_Sorter100|15742_ ,
    \new_Sorter100|15743_ , \new_Sorter100|15744_ , \new_Sorter100|15745_ ,
    \new_Sorter100|15746_ , \new_Sorter100|15747_ , \new_Sorter100|15748_ ,
    \new_Sorter100|15749_ , \new_Sorter100|15750_ , \new_Sorter100|15751_ ,
    \new_Sorter100|15752_ , \new_Sorter100|15753_ , \new_Sorter100|15754_ ,
    \new_Sorter100|15755_ , \new_Sorter100|15756_ , \new_Sorter100|15757_ ,
    \new_Sorter100|15758_ , \new_Sorter100|15759_ , \new_Sorter100|15760_ ,
    \new_Sorter100|15761_ , \new_Sorter100|15762_ , \new_Sorter100|15763_ ,
    \new_Sorter100|15764_ , \new_Sorter100|15765_ , \new_Sorter100|15766_ ,
    \new_Sorter100|15767_ , \new_Sorter100|15768_ , \new_Sorter100|15769_ ,
    \new_Sorter100|15770_ , \new_Sorter100|15771_ , \new_Sorter100|15772_ ,
    \new_Sorter100|15773_ , \new_Sorter100|15774_ , \new_Sorter100|15775_ ,
    \new_Sorter100|15776_ , \new_Sorter100|15777_ , \new_Sorter100|15778_ ,
    \new_Sorter100|15779_ , \new_Sorter100|15780_ , \new_Sorter100|15781_ ,
    \new_Sorter100|15782_ , \new_Sorter100|15783_ , \new_Sorter100|15784_ ,
    \new_Sorter100|15785_ , \new_Sorter100|15786_ , \new_Sorter100|15787_ ,
    \new_Sorter100|15788_ , \new_Sorter100|15789_ , \new_Sorter100|15790_ ,
    \new_Sorter100|15791_ , \new_Sorter100|15792_ , \new_Sorter100|15793_ ,
    \new_Sorter100|15794_ , \new_Sorter100|15795_ , \new_Sorter100|15796_ ,
    \new_Sorter100|15797_ , \new_Sorter100|15798_ , \new_Sorter100|15800_ ,
    \new_Sorter100|15801_ , \new_Sorter100|15802_ , \new_Sorter100|15803_ ,
    \new_Sorter100|15804_ , \new_Sorter100|15805_ , \new_Sorter100|15806_ ,
    \new_Sorter100|15807_ , \new_Sorter100|15808_ , \new_Sorter100|15809_ ,
    \new_Sorter100|15810_ , \new_Sorter100|15811_ , \new_Sorter100|15812_ ,
    \new_Sorter100|15813_ , \new_Sorter100|15814_ , \new_Sorter100|15815_ ,
    \new_Sorter100|15816_ , \new_Sorter100|15817_ , \new_Sorter100|15818_ ,
    \new_Sorter100|15819_ , \new_Sorter100|15820_ , \new_Sorter100|15821_ ,
    \new_Sorter100|15822_ , \new_Sorter100|15823_ , \new_Sorter100|15824_ ,
    \new_Sorter100|15825_ , \new_Sorter100|15826_ , \new_Sorter100|15827_ ,
    \new_Sorter100|15828_ , \new_Sorter100|15829_ , \new_Sorter100|15830_ ,
    \new_Sorter100|15831_ , \new_Sorter100|15832_ , \new_Sorter100|15833_ ,
    \new_Sorter100|15834_ , \new_Sorter100|15835_ , \new_Sorter100|15836_ ,
    \new_Sorter100|15837_ , \new_Sorter100|15838_ , \new_Sorter100|15839_ ,
    \new_Sorter100|15840_ , \new_Sorter100|15841_ , \new_Sorter100|15842_ ,
    \new_Sorter100|15843_ , \new_Sorter100|15844_ , \new_Sorter100|15845_ ,
    \new_Sorter100|15846_ , \new_Sorter100|15847_ , \new_Sorter100|15848_ ,
    \new_Sorter100|15849_ , \new_Sorter100|15850_ , \new_Sorter100|15851_ ,
    \new_Sorter100|15852_ , \new_Sorter100|15853_ , \new_Sorter100|15854_ ,
    \new_Sorter100|15855_ , \new_Sorter100|15856_ , \new_Sorter100|15857_ ,
    \new_Sorter100|15858_ , \new_Sorter100|15859_ , \new_Sorter100|15860_ ,
    \new_Sorter100|15861_ , \new_Sorter100|15862_ , \new_Sorter100|15863_ ,
    \new_Sorter100|15864_ , \new_Sorter100|15865_ , \new_Sorter100|15866_ ,
    \new_Sorter100|15867_ , \new_Sorter100|15868_ , \new_Sorter100|15869_ ,
    \new_Sorter100|15870_ , \new_Sorter100|15871_ , \new_Sorter100|15872_ ,
    \new_Sorter100|15873_ , \new_Sorter100|15874_ , \new_Sorter100|15875_ ,
    \new_Sorter100|15876_ , \new_Sorter100|15877_ , \new_Sorter100|15878_ ,
    \new_Sorter100|15879_ , \new_Sorter100|15880_ , \new_Sorter100|15881_ ,
    \new_Sorter100|15882_ , \new_Sorter100|15883_ , \new_Sorter100|15884_ ,
    \new_Sorter100|15885_ , \new_Sorter100|15886_ , \new_Sorter100|15887_ ,
    \new_Sorter100|15888_ , \new_Sorter100|15889_ , \new_Sorter100|15890_ ,
    \new_Sorter100|15891_ , \new_Sorter100|15892_ , \new_Sorter100|15893_ ,
    \new_Sorter100|15894_ , \new_Sorter100|15895_ , \new_Sorter100|15896_ ,
    \new_Sorter100|15897_ , \new_Sorter100|15898_ , \new_Sorter100|15899_ ,
    \new_Sorter100|15900_ , \new_Sorter100|15999_ , \new_Sorter100|15901_ ,
    \new_Sorter100|15902_ , \new_Sorter100|15903_ , \new_Sorter100|15904_ ,
    \new_Sorter100|15905_ , \new_Sorter100|15906_ , \new_Sorter100|15907_ ,
    \new_Sorter100|15908_ , \new_Sorter100|15909_ , \new_Sorter100|15910_ ,
    \new_Sorter100|15911_ , \new_Sorter100|15912_ , \new_Sorter100|15913_ ,
    \new_Sorter100|15914_ , \new_Sorter100|15915_ , \new_Sorter100|15916_ ,
    \new_Sorter100|15917_ , \new_Sorter100|15918_ , \new_Sorter100|15919_ ,
    \new_Sorter100|15920_ , \new_Sorter100|15921_ , \new_Sorter100|15922_ ,
    \new_Sorter100|15923_ , \new_Sorter100|15924_ , \new_Sorter100|15925_ ,
    \new_Sorter100|15926_ , \new_Sorter100|15927_ , \new_Sorter100|15928_ ,
    \new_Sorter100|15929_ , \new_Sorter100|15930_ , \new_Sorter100|15931_ ,
    \new_Sorter100|15932_ , \new_Sorter100|15933_ , \new_Sorter100|15934_ ,
    \new_Sorter100|15935_ , \new_Sorter100|15936_ , \new_Sorter100|15937_ ,
    \new_Sorter100|15938_ , \new_Sorter100|15939_ , \new_Sorter100|15940_ ,
    \new_Sorter100|15941_ , \new_Sorter100|15942_ , \new_Sorter100|15943_ ,
    \new_Sorter100|15944_ , \new_Sorter100|15945_ , \new_Sorter100|15946_ ,
    \new_Sorter100|15947_ , \new_Sorter100|15948_ , \new_Sorter100|15949_ ,
    \new_Sorter100|15950_ , \new_Sorter100|15951_ , \new_Sorter100|15952_ ,
    \new_Sorter100|15953_ , \new_Sorter100|15954_ , \new_Sorter100|15955_ ,
    \new_Sorter100|15956_ , \new_Sorter100|15957_ , \new_Sorter100|15958_ ,
    \new_Sorter100|15959_ , \new_Sorter100|15960_ , \new_Sorter100|15961_ ,
    \new_Sorter100|15962_ , \new_Sorter100|15963_ , \new_Sorter100|15964_ ,
    \new_Sorter100|15965_ , \new_Sorter100|15966_ , \new_Sorter100|15967_ ,
    \new_Sorter100|15968_ , \new_Sorter100|15969_ , \new_Sorter100|15970_ ,
    \new_Sorter100|15971_ , \new_Sorter100|15972_ , \new_Sorter100|15973_ ,
    \new_Sorter100|15974_ , \new_Sorter100|15975_ , \new_Sorter100|15976_ ,
    \new_Sorter100|15977_ , \new_Sorter100|15978_ , \new_Sorter100|15979_ ,
    \new_Sorter100|15980_ , \new_Sorter100|15981_ , \new_Sorter100|15982_ ,
    \new_Sorter100|15983_ , \new_Sorter100|15984_ , \new_Sorter100|15985_ ,
    \new_Sorter100|15986_ , \new_Sorter100|15987_ , \new_Sorter100|15988_ ,
    \new_Sorter100|15989_ , \new_Sorter100|15990_ , \new_Sorter100|15991_ ,
    \new_Sorter100|15992_ , \new_Sorter100|15993_ , \new_Sorter100|15994_ ,
    \new_Sorter100|15995_ , \new_Sorter100|15996_ , \new_Sorter100|15997_ ,
    \new_Sorter100|15998_ , \new_Sorter100|16000_ , \new_Sorter100|16001_ ,
    \new_Sorter100|16002_ , \new_Sorter100|16003_ , \new_Sorter100|16004_ ,
    \new_Sorter100|16005_ , \new_Sorter100|16006_ , \new_Sorter100|16007_ ,
    \new_Sorter100|16008_ , \new_Sorter100|16009_ , \new_Sorter100|16010_ ,
    \new_Sorter100|16011_ , \new_Sorter100|16012_ , \new_Sorter100|16013_ ,
    \new_Sorter100|16014_ , \new_Sorter100|16015_ , \new_Sorter100|16016_ ,
    \new_Sorter100|16017_ , \new_Sorter100|16018_ , \new_Sorter100|16019_ ,
    \new_Sorter100|16020_ , \new_Sorter100|16021_ , \new_Sorter100|16022_ ,
    \new_Sorter100|16023_ , \new_Sorter100|16024_ , \new_Sorter100|16025_ ,
    \new_Sorter100|16026_ , \new_Sorter100|16027_ , \new_Sorter100|16028_ ,
    \new_Sorter100|16029_ , \new_Sorter100|16030_ , \new_Sorter100|16031_ ,
    \new_Sorter100|16032_ , \new_Sorter100|16033_ , \new_Sorter100|16034_ ,
    \new_Sorter100|16035_ , \new_Sorter100|16036_ , \new_Sorter100|16037_ ,
    \new_Sorter100|16038_ , \new_Sorter100|16039_ , \new_Sorter100|16040_ ,
    \new_Sorter100|16041_ , \new_Sorter100|16042_ , \new_Sorter100|16043_ ,
    \new_Sorter100|16044_ , \new_Sorter100|16045_ , \new_Sorter100|16046_ ,
    \new_Sorter100|16047_ , \new_Sorter100|16048_ , \new_Sorter100|16049_ ,
    \new_Sorter100|16050_ , \new_Sorter100|16051_ , \new_Sorter100|16052_ ,
    \new_Sorter100|16053_ , \new_Sorter100|16054_ , \new_Sorter100|16055_ ,
    \new_Sorter100|16056_ , \new_Sorter100|16057_ , \new_Sorter100|16058_ ,
    \new_Sorter100|16059_ , \new_Sorter100|16060_ , \new_Sorter100|16061_ ,
    \new_Sorter100|16062_ , \new_Sorter100|16063_ , \new_Sorter100|16064_ ,
    \new_Sorter100|16065_ , \new_Sorter100|16066_ , \new_Sorter100|16067_ ,
    \new_Sorter100|16068_ , \new_Sorter100|16069_ , \new_Sorter100|16070_ ,
    \new_Sorter100|16071_ , \new_Sorter100|16072_ , \new_Sorter100|16073_ ,
    \new_Sorter100|16074_ , \new_Sorter100|16075_ , \new_Sorter100|16076_ ,
    \new_Sorter100|16077_ , \new_Sorter100|16078_ , \new_Sorter100|16079_ ,
    \new_Sorter100|16080_ , \new_Sorter100|16081_ , \new_Sorter100|16082_ ,
    \new_Sorter100|16083_ , \new_Sorter100|16084_ , \new_Sorter100|16085_ ,
    \new_Sorter100|16086_ , \new_Sorter100|16087_ , \new_Sorter100|16088_ ,
    \new_Sorter100|16089_ , \new_Sorter100|16090_ , \new_Sorter100|16091_ ,
    \new_Sorter100|16092_ , \new_Sorter100|16093_ , \new_Sorter100|16094_ ,
    \new_Sorter100|16095_ , \new_Sorter100|16096_ , \new_Sorter100|16097_ ,
    \new_Sorter100|16098_ , \new_Sorter100|16099_ , \new_Sorter100|16100_ ,
    \new_Sorter100|16199_ , \new_Sorter100|16101_ , \new_Sorter100|16102_ ,
    \new_Sorter100|16103_ , \new_Sorter100|16104_ , \new_Sorter100|16105_ ,
    \new_Sorter100|16106_ , \new_Sorter100|16107_ , \new_Sorter100|16108_ ,
    \new_Sorter100|16109_ , \new_Sorter100|16110_ , \new_Sorter100|16111_ ,
    \new_Sorter100|16112_ , \new_Sorter100|16113_ , \new_Sorter100|16114_ ,
    \new_Sorter100|16115_ , \new_Sorter100|16116_ , \new_Sorter100|16117_ ,
    \new_Sorter100|16118_ , \new_Sorter100|16119_ , \new_Sorter100|16120_ ,
    \new_Sorter100|16121_ , \new_Sorter100|16122_ , \new_Sorter100|16123_ ,
    \new_Sorter100|16124_ , \new_Sorter100|16125_ , \new_Sorter100|16126_ ,
    \new_Sorter100|16127_ , \new_Sorter100|16128_ , \new_Sorter100|16129_ ,
    \new_Sorter100|16130_ , \new_Sorter100|16131_ , \new_Sorter100|16132_ ,
    \new_Sorter100|16133_ , \new_Sorter100|16134_ , \new_Sorter100|16135_ ,
    \new_Sorter100|16136_ , \new_Sorter100|16137_ , \new_Sorter100|16138_ ,
    \new_Sorter100|16139_ , \new_Sorter100|16140_ , \new_Sorter100|16141_ ,
    \new_Sorter100|16142_ , \new_Sorter100|16143_ , \new_Sorter100|16144_ ,
    \new_Sorter100|16145_ , \new_Sorter100|16146_ , \new_Sorter100|16147_ ,
    \new_Sorter100|16148_ , \new_Sorter100|16149_ , \new_Sorter100|16150_ ,
    \new_Sorter100|16151_ , \new_Sorter100|16152_ , \new_Sorter100|16153_ ,
    \new_Sorter100|16154_ , \new_Sorter100|16155_ , \new_Sorter100|16156_ ,
    \new_Sorter100|16157_ , \new_Sorter100|16158_ , \new_Sorter100|16159_ ,
    \new_Sorter100|16160_ , \new_Sorter100|16161_ , \new_Sorter100|16162_ ,
    \new_Sorter100|16163_ , \new_Sorter100|16164_ , \new_Sorter100|16165_ ,
    \new_Sorter100|16166_ , \new_Sorter100|16167_ , \new_Sorter100|16168_ ,
    \new_Sorter100|16169_ , \new_Sorter100|16170_ , \new_Sorter100|16171_ ,
    \new_Sorter100|16172_ , \new_Sorter100|16173_ , \new_Sorter100|16174_ ,
    \new_Sorter100|16175_ , \new_Sorter100|16176_ , \new_Sorter100|16177_ ,
    \new_Sorter100|16178_ , \new_Sorter100|16179_ , \new_Sorter100|16180_ ,
    \new_Sorter100|16181_ , \new_Sorter100|16182_ , \new_Sorter100|16183_ ,
    \new_Sorter100|16184_ , \new_Sorter100|16185_ , \new_Sorter100|16186_ ,
    \new_Sorter100|16187_ , \new_Sorter100|16188_ , \new_Sorter100|16189_ ,
    \new_Sorter100|16190_ , \new_Sorter100|16191_ , \new_Sorter100|16192_ ,
    \new_Sorter100|16193_ , \new_Sorter100|16194_ , \new_Sorter100|16195_ ,
    \new_Sorter100|16196_ , \new_Sorter100|16197_ , \new_Sorter100|16198_ ,
    \new_Sorter100|16200_ , \new_Sorter100|16201_ , \new_Sorter100|16202_ ,
    \new_Sorter100|16203_ , \new_Sorter100|16204_ , \new_Sorter100|16205_ ,
    \new_Sorter100|16206_ , \new_Sorter100|16207_ , \new_Sorter100|16208_ ,
    \new_Sorter100|16209_ , \new_Sorter100|16210_ , \new_Sorter100|16211_ ,
    \new_Sorter100|16212_ , \new_Sorter100|16213_ , \new_Sorter100|16214_ ,
    \new_Sorter100|16215_ , \new_Sorter100|16216_ , \new_Sorter100|16217_ ,
    \new_Sorter100|16218_ , \new_Sorter100|16219_ , \new_Sorter100|16220_ ,
    \new_Sorter100|16221_ , \new_Sorter100|16222_ , \new_Sorter100|16223_ ,
    \new_Sorter100|16224_ , \new_Sorter100|16225_ , \new_Sorter100|16226_ ,
    \new_Sorter100|16227_ , \new_Sorter100|16228_ , \new_Sorter100|16229_ ,
    \new_Sorter100|16230_ , \new_Sorter100|16231_ , \new_Sorter100|16232_ ,
    \new_Sorter100|16233_ , \new_Sorter100|16234_ , \new_Sorter100|16235_ ,
    \new_Sorter100|16236_ , \new_Sorter100|16237_ , \new_Sorter100|16238_ ,
    \new_Sorter100|16239_ , \new_Sorter100|16240_ , \new_Sorter100|16241_ ,
    \new_Sorter100|16242_ , \new_Sorter100|16243_ , \new_Sorter100|16244_ ,
    \new_Sorter100|16245_ , \new_Sorter100|16246_ , \new_Sorter100|16247_ ,
    \new_Sorter100|16248_ , \new_Sorter100|16249_ , \new_Sorter100|16250_ ,
    \new_Sorter100|16251_ , \new_Sorter100|16252_ , \new_Sorter100|16253_ ,
    \new_Sorter100|16254_ , \new_Sorter100|16255_ , \new_Sorter100|16256_ ,
    \new_Sorter100|16257_ , \new_Sorter100|16258_ , \new_Sorter100|16259_ ,
    \new_Sorter100|16260_ , \new_Sorter100|16261_ , \new_Sorter100|16262_ ,
    \new_Sorter100|16263_ , \new_Sorter100|16264_ , \new_Sorter100|16265_ ,
    \new_Sorter100|16266_ , \new_Sorter100|16267_ , \new_Sorter100|16268_ ,
    \new_Sorter100|16269_ , \new_Sorter100|16270_ , \new_Sorter100|16271_ ,
    \new_Sorter100|16272_ , \new_Sorter100|16273_ , \new_Sorter100|16274_ ,
    \new_Sorter100|16275_ , \new_Sorter100|16276_ , \new_Sorter100|16277_ ,
    \new_Sorter100|16278_ , \new_Sorter100|16279_ , \new_Sorter100|16280_ ,
    \new_Sorter100|16281_ , \new_Sorter100|16282_ , \new_Sorter100|16283_ ,
    \new_Sorter100|16284_ , \new_Sorter100|16285_ , \new_Sorter100|16286_ ,
    \new_Sorter100|16287_ , \new_Sorter100|16288_ , \new_Sorter100|16289_ ,
    \new_Sorter100|16290_ , \new_Sorter100|16291_ , \new_Sorter100|16292_ ,
    \new_Sorter100|16293_ , \new_Sorter100|16294_ , \new_Sorter100|16295_ ,
    \new_Sorter100|16296_ , \new_Sorter100|16297_ , \new_Sorter100|16298_ ,
    \new_Sorter100|16299_ , \new_Sorter100|16300_ , \new_Sorter100|16399_ ,
    \new_Sorter100|16301_ , \new_Sorter100|16302_ , \new_Sorter100|16303_ ,
    \new_Sorter100|16304_ , \new_Sorter100|16305_ , \new_Sorter100|16306_ ,
    \new_Sorter100|16307_ , \new_Sorter100|16308_ , \new_Sorter100|16309_ ,
    \new_Sorter100|16310_ , \new_Sorter100|16311_ , \new_Sorter100|16312_ ,
    \new_Sorter100|16313_ , \new_Sorter100|16314_ , \new_Sorter100|16315_ ,
    \new_Sorter100|16316_ , \new_Sorter100|16317_ , \new_Sorter100|16318_ ,
    \new_Sorter100|16319_ , \new_Sorter100|16320_ , \new_Sorter100|16321_ ,
    \new_Sorter100|16322_ , \new_Sorter100|16323_ , \new_Sorter100|16324_ ,
    \new_Sorter100|16325_ , \new_Sorter100|16326_ , \new_Sorter100|16327_ ,
    \new_Sorter100|16328_ , \new_Sorter100|16329_ , \new_Sorter100|16330_ ,
    \new_Sorter100|16331_ , \new_Sorter100|16332_ , \new_Sorter100|16333_ ,
    \new_Sorter100|16334_ , \new_Sorter100|16335_ , \new_Sorter100|16336_ ,
    \new_Sorter100|16337_ , \new_Sorter100|16338_ , \new_Sorter100|16339_ ,
    \new_Sorter100|16340_ , \new_Sorter100|16341_ , \new_Sorter100|16342_ ,
    \new_Sorter100|16343_ , \new_Sorter100|16344_ , \new_Sorter100|16345_ ,
    \new_Sorter100|16346_ , \new_Sorter100|16347_ , \new_Sorter100|16348_ ,
    \new_Sorter100|16349_ , \new_Sorter100|16350_ , \new_Sorter100|16351_ ,
    \new_Sorter100|16352_ , \new_Sorter100|16353_ , \new_Sorter100|16354_ ,
    \new_Sorter100|16355_ , \new_Sorter100|16356_ , \new_Sorter100|16357_ ,
    \new_Sorter100|16358_ , \new_Sorter100|16359_ , \new_Sorter100|16360_ ,
    \new_Sorter100|16361_ , \new_Sorter100|16362_ , \new_Sorter100|16363_ ,
    \new_Sorter100|16364_ , \new_Sorter100|16365_ , \new_Sorter100|16366_ ,
    \new_Sorter100|16367_ , \new_Sorter100|16368_ , \new_Sorter100|16369_ ,
    \new_Sorter100|16370_ , \new_Sorter100|16371_ , \new_Sorter100|16372_ ,
    \new_Sorter100|16373_ , \new_Sorter100|16374_ , \new_Sorter100|16375_ ,
    \new_Sorter100|16376_ , \new_Sorter100|16377_ , \new_Sorter100|16378_ ,
    \new_Sorter100|16379_ , \new_Sorter100|16380_ , \new_Sorter100|16381_ ,
    \new_Sorter100|16382_ , \new_Sorter100|16383_ , \new_Sorter100|16384_ ,
    \new_Sorter100|16385_ , \new_Sorter100|16386_ , \new_Sorter100|16387_ ,
    \new_Sorter100|16388_ , \new_Sorter100|16389_ , \new_Sorter100|16390_ ,
    \new_Sorter100|16391_ , \new_Sorter100|16392_ , \new_Sorter100|16393_ ,
    \new_Sorter100|16394_ , \new_Sorter100|16395_ , \new_Sorter100|16396_ ,
    \new_Sorter100|16397_ , \new_Sorter100|16398_ , \new_Sorter100|16400_ ,
    \new_Sorter100|16401_ , \new_Sorter100|16402_ , \new_Sorter100|16403_ ,
    \new_Sorter100|16404_ , \new_Sorter100|16405_ , \new_Sorter100|16406_ ,
    \new_Sorter100|16407_ , \new_Sorter100|16408_ , \new_Sorter100|16409_ ,
    \new_Sorter100|16410_ , \new_Sorter100|16411_ , \new_Sorter100|16412_ ,
    \new_Sorter100|16413_ , \new_Sorter100|16414_ , \new_Sorter100|16415_ ,
    \new_Sorter100|16416_ , \new_Sorter100|16417_ , \new_Sorter100|16418_ ,
    \new_Sorter100|16419_ , \new_Sorter100|16420_ , \new_Sorter100|16421_ ,
    \new_Sorter100|16422_ , \new_Sorter100|16423_ , \new_Sorter100|16424_ ,
    \new_Sorter100|16425_ , \new_Sorter100|16426_ , \new_Sorter100|16427_ ,
    \new_Sorter100|16428_ , \new_Sorter100|16429_ , \new_Sorter100|16430_ ,
    \new_Sorter100|16431_ , \new_Sorter100|16432_ , \new_Sorter100|16433_ ,
    \new_Sorter100|16434_ , \new_Sorter100|16435_ , \new_Sorter100|16436_ ,
    \new_Sorter100|16437_ , \new_Sorter100|16438_ , \new_Sorter100|16439_ ,
    \new_Sorter100|16440_ , \new_Sorter100|16441_ , \new_Sorter100|16442_ ,
    \new_Sorter100|16443_ , \new_Sorter100|16444_ , \new_Sorter100|16445_ ,
    \new_Sorter100|16446_ , \new_Sorter100|16447_ , \new_Sorter100|16448_ ,
    \new_Sorter100|16449_ , \new_Sorter100|16450_ , \new_Sorter100|16451_ ,
    \new_Sorter100|16452_ , \new_Sorter100|16453_ , \new_Sorter100|16454_ ,
    \new_Sorter100|16455_ , \new_Sorter100|16456_ , \new_Sorter100|16457_ ,
    \new_Sorter100|16458_ , \new_Sorter100|16459_ , \new_Sorter100|16460_ ,
    \new_Sorter100|16461_ , \new_Sorter100|16462_ , \new_Sorter100|16463_ ,
    \new_Sorter100|16464_ , \new_Sorter100|16465_ , \new_Sorter100|16466_ ,
    \new_Sorter100|16467_ , \new_Sorter100|16468_ , \new_Sorter100|16469_ ,
    \new_Sorter100|16470_ , \new_Sorter100|16471_ , \new_Sorter100|16472_ ,
    \new_Sorter100|16473_ , \new_Sorter100|16474_ , \new_Sorter100|16475_ ,
    \new_Sorter100|16476_ , \new_Sorter100|16477_ , \new_Sorter100|16478_ ,
    \new_Sorter100|16479_ , \new_Sorter100|16480_ , \new_Sorter100|16481_ ,
    \new_Sorter100|16482_ , \new_Sorter100|16483_ , \new_Sorter100|16484_ ,
    \new_Sorter100|16485_ , \new_Sorter100|16486_ , \new_Sorter100|16487_ ,
    \new_Sorter100|16488_ , \new_Sorter100|16489_ , \new_Sorter100|16490_ ,
    \new_Sorter100|16491_ , \new_Sorter100|16492_ , \new_Sorter100|16493_ ,
    \new_Sorter100|16494_ , \new_Sorter100|16495_ , \new_Sorter100|16496_ ,
    \new_Sorter100|16497_ , \new_Sorter100|16498_ , \new_Sorter100|16499_ ,
    \new_Sorter100|16500_ , \new_Sorter100|16599_ , \new_Sorter100|16501_ ,
    \new_Sorter100|16502_ , \new_Sorter100|16503_ , \new_Sorter100|16504_ ,
    \new_Sorter100|16505_ , \new_Sorter100|16506_ , \new_Sorter100|16507_ ,
    \new_Sorter100|16508_ , \new_Sorter100|16509_ , \new_Sorter100|16510_ ,
    \new_Sorter100|16511_ , \new_Sorter100|16512_ , \new_Sorter100|16513_ ,
    \new_Sorter100|16514_ , \new_Sorter100|16515_ , \new_Sorter100|16516_ ,
    \new_Sorter100|16517_ , \new_Sorter100|16518_ , \new_Sorter100|16519_ ,
    \new_Sorter100|16520_ , \new_Sorter100|16521_ , \new_Sorter100|16522_ ,
    \new_Sorter100|16523_ , \new_Sorter100|16524_ , \new_Sorter100|16525_ ,
    \new_Sorter100|16526_ , \new_Sorter100|16527_ , \new_Sorter100|16528_ ,
    \new_Sorter100|16529_ , \new_Sorter100|16530_ , \new_Sorter100|16531_ ,
    \new_Sorter100|16532_ , \new_Sorter100|16533_ , \new_Sorter100|16534_ ,
    \new_Sorter100|16535_ , \new_Sorter100|16536_ , \new_Sorter100|16537_ ,
    \new_Sorter100|16538_ , \new_Sorter100|16539_ , \new_Sorter100|16540_ ,
    \new_Sorter100|16541_ , \new_Sorter100|16542_ , \new_Sorter100|16543_ ,
    \new_Sorter100|16544_ , \new_Sorter100|16545_ , \new_Sorter100|16546_ ,
    \new_Sorter100|16547_ , \new_Sorter100|16548_ , \new_Sorter100|16549_ ,
    \new_Sorter100|16550_ , \new_Sorter100|16551_ , \new_Sorter100|16552_ ,
    \new_Sorter100|16553_ , \new_Sorter100|16554_ , \new_Sorter100|16555_ ,
    \new_Sorter100|16556_ , \new_Sorter100|16557_ , \new_Sorter100|16558_ ,
    \new_Sorter100|16559_ , \new_Sorter100|16560_ , \new_Sorter100|16561_ ,
    \new_Sorter100|16562_ , \new_Sorter100|16563_ , \new_Sorter100|16564_ ,
    \new_Sorter100|16565_ , \new_Sorter100|16566_ , \new_Sorter100|16567_ ,
    \new_Sorter100|16568_ , \new_Sorter100|16569_ , \new_Sorter100|16570_ ,
    \new_Sorter100|16571_ , \new_Sorter100|16572_ , \new_Sorter100|16573_ ,
    \new_Sorter100|16574_ , \new_Sorter100|16575_ , \new_Sorter100|16576_ ,
    \new_Sorter100|16577_ , \new_Sorter100|16578_ , \new_Sorter100|16579_ ,
    \new_Sorter100|16580_ , \new_Sorter100|16581_ , \new_Sorter100|16582_ ,
    \new_Sorter100|16583_ , \new_Sorter100|16584_ , \new_Sorter100|16585_ ,
    \new_Sorter100|16586_ , \new_Sorter100|16587_ , \new_Sorter100|16588_ ,
    \new_Sorter100|16589_ , \new_Sorter100|16590_ , \new_Sorter100|16591_ ,
    \new_Sorter100|16592_ , \new_Sorter100|16593_ , \new_Sorter100|16594_ ,
    \new_Sorter100|16595_ , \new_Sorter100|16596_ , \new_Sorter100|16597_ ,
    \new_Sorter100|16598_ , \new_Sorter100|16600_ , \new_Sorter100|16601_ ,
    \new_Sorter100|16602_ , \new_Sorter100|16603_ , \new_Sorter100|16604_ ,
    \new_Sorter100|16605_ , \new_Sorter100|16606_ , \new_Sorter100|16607_ ,
    \new_Sorter100|16608_ , \new_Sorter100|16609_ , \new_Sorter100|16610_ ,
    \new_Sorter100|16611_ , \new_Sorter100|16612_ , \new_Sorter100|16613_ ,
    \new_Sorter100|16614_ , \new_Sorter100|16615_ , \new_Sorter100|16616_ ,
    \new_Sorter100|16617_ , \new_Sorter100|16618_ , \new_Sorter100|16619_ ,
    \new_Sorter100|16620_ , \new_Sorter100|16621_ , \new_Sorter100|16622_ ,
    \new_Sorter100|16623_ , \new_Sorter100|16624_ , \new_Sorter100|16625_ ,
    \new_Sorter100|16626_ , \new_Sorter100|16627_ , \new_Sorter100|16628_ ,
    \new_Sorter100|16629_ , \new_Sorter100|16630_ , \new_Sorter100|16631_ ,
    \new_Sorter100|16632_ , \new_Sorter100|16633_ , \new_Sorter100|16634_ ,
    \new_Sorter100|16635_ , \new_Sorter100|16636_ , \new_Sorter100|16637_ ,
    \new_Sorter100|16638_ , \new_Sorter100|16639_ , \new_Sorter100|16640_ ,
    \new_Sorter100|16641_ , \new_Sorter100|16642_ , \new_Sorter100|16643_ ,
    \new_Sorter100|16644_ , \new_Sorter100|16645_ , \new_Sorter100|16646_ ,
    \new_Sorter100|16647_ , \new_Sorter100|16648_ , \new_Sorter100|16649_ ,
    \new_Sorter100|16650_ , \new_Sorter100|16651_ , \new_Sorter100|16652_ ,
    \new_Sorter100|16653_ , \new_Sorter100|16654_ , \new_Sorter100|16655_ ,
    \new_Sorter100|16656_ , \new_Sorter100|16657_ , \new_Sorter100|16658_ ,
    \new_Sorter100|16659_ , \new_Sorter100|16660_ , \new_Sorter100|16661_ ,
    \new_Sorter100|16662_ , \new_Sorter100|16663_ , \new_Sorter100|16664_ ,
    \new_Sorter100|16665_ , \new_Sorter100|16666_ , \new_Sorter100|16667_ ,
    \new_Sorter100|16668_ , \new_Sorter100|16669_ , \new_Sorter100|16670_ ,
    \new_Sorter100|16671_ , \new_Sorter100|16672_ , \new_Sorter100|16673_ ,
    \new_Sorter100|16674_ , \new_Sorter100|16675_ , \new_Sorter100|16676_ ,
    \new_Sorter100|16677_ , \new_Sorter100|16678_ , \new_Sorter100|16679_ ,
    \new_Sorter100|16680_ , \new_Sorter100|16681_ , \new_Sorter100|16682_ ,
    \new_Sorter100|16683_ , \new_Sorter100|16684_ , \new_Sorter100|16685_ ,
    \new_Sorter100|16686_ , \new_Sorter100|16687_ , \new_Sorter100|16688_ ,
    \new_Sorter100|16689_ , \new_Sorter100|16690_ , \new_Sorter100|16691_ ,
    \new_Sorter100|16692_ , \new_Sorter100|16693_ , \new_Sorter100|16694_ ,
    \new_Sorter100|16695_ , \new_Sorter100|16696_ , \new_Sorter100|16697_ ,
    \new_Sorter100|16698_ , \new_Sorter100|16699_ , \new_Sorter100|16700_ ,
    \new_Sorter100|16799_ , \new_Sorter100|16701_ , \new_Sorter100|16702_ ,
    \new_Sorter100|16703_ , \new_Sorter100|16704_ , \new_Sorter100|16705_ ,
    \new_Sorter100|16706_ , \new_Sorter100|16707_ , \new_Sorter100|16708_ ,
    \new_Sorter100|16709_ , \new_Sorter100|16710_ , \new_Sorter100|16711_ ,
    \new_Sorter100|16712_ , \new_Sorter100|16713_ , \new_Sorter100|16714_ ,
    \new_Sorter100|16715_ , \new_Sorter100|16716_ , \new_Sorter100|16717_ ,
    \new_Sorter100|16718_ , \new_Sorter100|16719_ , \new_Sorter100|16720_ ,
    \new_Sorter100|16721_ , \new_Sorter100|16722_ , \new_Sorter100|16723_ ,
    \new_Sorter100|16724_ , \new_Sorter100|16725_ , \new_Sorter100|16726_ ,
    \new_Sorter100|16727_ , \new_Sorter100|16728_ , \new_Sorter100|16729_ ,
    \new_Sorter100|16730_ , \new_Sorter100|16731_ , \new_Sorter100|16732_ ,
    \new_Sorter100|16733_ , \new_Sorter100|16734_ , \new_Sorter100|16735_ ,
    \new_Sorter100|16736_ , \new_Sorter100|16737_ , \new_Sorter100|16738_ ,
    \new_Sorter100|16739_ , \new_Sorter100|16740_ , \new_Sorter100|16741_ ,
    \new_Sorter100|16742_ , \new_Sorter100|16743_ , \new_Sorter100|16744_ ,
    \new_Sorter100|16745_ , \new_Sorter100|16746_ , \new_Sorter100|16747_ ,
    \new_Sorter100|16748_ , \new_Sorter100|16749_ , \new_Sorter100|16750_ ,
    \new_Sorter100|16751_ , \new_Sorter100|16752_ , \new_Sorter100|16753_ ,
    \new_Sorter100|16754_ , \new_Sorter100|16755_ , \new_Sorter100|16756_ ,
    \new_Sorter100|16757_ , \new_Sorter100|16758_ , \new_Sorter100|16759_ ,
    \new_Sorter100|16760_ , \new_Sorter100|16761_ , \new_Sorter100|16762_ ,
    \new_Sorter100|16763_ , \new_Sorter100|16764_ , \new_Sorter100|16765_ ,
    \new_Sorter100|16766_ , \new_Sorter100|16767_ , \new_Sorter100|16768_ ,
    \new_Sorter100|16769_ , \new_Sorter100|16770_ , \new_Sorter100|16771_ ,
    \new_Sorter100|16772_ , \new_Sorter100|16773_ , \new_Sorter100|16774_ ,
    \new_Sorter100|16775_ , \new_Sorter100|16776_ , \new_Sorter100|16777_ ,
    \new_Sorter100|16778_ , \new_Sorter100|16779_ , \new_Sorter100|16780_ ,
    \new_Sorter100|16781_ , \new_Sorter100|16782_ , \new_Sorter100|16783_ ,
    \new_Sorter100|16784_ , \new_Sorter100|16785_ , \new_Sorter100|16786_ ,
    \new_Sorter100|16787_ , \new_Sorter100|16788_ , \new_Sorter100|16789_ ,
    \new_Sorter100|16790_ , \new_Sorter100|16791_ , \new_Sorter100|16792_ ,
    \new_Sorter100|16793_ , \new_Sorter100|16794_ , \new_Sorter100|16795_ ,
    \new_Sorter100|16796_ , \new_Sorter100|16797_ , \new_Sorter100|16798_ ,
    \new_Sorter100|16800_ , \new_Sorter100|16801_ , \new_Sorter100|16802_ ,
    \new_Sorter100|16803_ , \new_Sorter100|16804_ , \new_Sorter100|16805_ ,
    \new_Sorter100|16806_ , \new_Sorter100|16807_ , \new_Sorter100|16808_ ,
    \new_Sorter100|16809_ , \new_Sorter100|16810_ , \new_Sorter100|16811_ ,
    \new_Sorter100|16812_ , \new_Sorter100|16813_ , \new_Sorter100|16814_ ,
    \new_Sorter100|16815_ , \new_Sorter100|16816_ , \new_Sorter100|16817_ ,
    \new_Sorter100|16818_ , \new_Sorter100|16819_ , \new_Sorter100|16820_ ,
    \new_Sorter100|16821_ , \new_Sorter100|16822_ , \new_Sorter100|16823_ ,
    \new_Sorter100|16824_ , \new_Sorter100|16825_ , \new_Sorter100|16826_ ,
    \new_Sorter100|16827_ , \new_Sorter100|16828_ , \new_Sorter100|16829_ ,
    \new_Sorter100|16830_ , \new_Sorter100|16831_ , \new_Sorter100|16832_ ,
    \new_Sorter100|16833_ , \new_Sorter100|16834_ , \new_Sorter100|16835_ ,
    \new_Sorter100|16836_ , \new_Sorter100|16837_ , \new_Sorter100|16838_ ,
    \new_Sorter100|16839_ , \new_Sorter100|16840_ , \new_Sorter100|16841_ ,
    \new_Sorter100|16842_ , \new_Sorter100|16843_ , \new_Sorter100|16844_ ,
    \new_Sorter100|16845_ , \new_Sorter100|16846_ , \new_Sorter100|16847_ ,
    \new_Sorter100|16848_ , \new_Sorter100|16849_ , \new_Sorter100|16850_ ,
    \new_Sorter100|16851_ , \new_Sorter100|16852_ , \new_Sorter100|16853_ ,
    \new_Sorter100|16854_ , \new_Sorter100|16855_ , \new_Sorter100|16856_ ,
    \new_Sorter100|16857_ , \new_Sorter100|16858_ , \new_Sorter100|16859_ ,
    \new_Sorter100|16860_ , \new_Sorter100|16861_ , \new_Sorter100|16862_ ,
    \new_Sorter100|16863_ , \new_Sorter100|16864_ , \new_Sorter100|16865_ ,
    \new_Sorter100|16866_ , \new_Sorter100|16867_ , \new_Sorter100|16868_ ,
    \new_Sorter100|16869_ , \new_Sorter100|16870_ , \new_Sorter100|16871_ ,
    \new_Sorter100|16872_ , \new_Sorter100|16873_ , \new_Sorter100|16874_ ,
    \new_Sorter100|16875_ , \new_Sorter100|16876_ , \new_Sorter100|16877_ ,
    \new_Sorter100|16878_ , \new_Sorter100|16879_ , \new_Sorter100|16880_ ,
    \new_Sorter100|16881_ , \new_Sorter100|16882_ , \new_Sorter100|16883_ ,
    \new_Sorter100|16884_ , \new_Sorter100|16885_ , \new_Sorter100|16886_ ,
    \new_Sorter100|16887_ , \new_Sorter100|16888_ , \new_Sorter100|16889_ ,
    \new_Sorter100|16890_ , \new_Sorter100|16891_ , \new_Sorter100|16892_ ,
    \new_Sorter100|16893_ , \new_Sorter100|16894_ , \new_Sorter100|16895_ ,
    \new_Sorter100|16896_ , \new_Sorter100|16897_ , \new_Sorter100|16898_ ,
    \new_Sorter100|16899_ , \new_Sorter100|16900_ , \new_Sorter100|16999_ ,
    \new_Sorter100|16901_ , \new_Sorter100|16902_ , \new_Sorter100|16903_ ,
    \new_Sorter100|16904_ , \new_Sorter100|16905_ , \new_Sorter100|16906_ ,
    \new_Sorter100|16907_ , \new_Sorter100|16908_ , \new_Sorter100|16909_ ,
    \new_Sorter100|16910_ , \new_Sorter100|16911_ , \new_Sorter100|16912_ ,
    \new_Sorter100|16913_ , \new_Sorter100|16914_ , \new_Sorter100|16915_ ,
    \new_Sorter100|16916_ , \new_Sorter100|16917_ , \new_Sorter100|16918_ ,
    \new_Sorter100|16919_ , \new_Sorter100|16920_ , \new_Sorter100|16921_ ,
    \new_Sorter100|16922_ , \new_Sorter100|16923_ , \new_Sorter100|16924_ ,
    \new_Sorter100|16925_ , \new_Sorter100|16926_ , \new_Sorter100|16927_ ,
    \new_Sorter100|16928_ , \new_Sorter100|16929_ , \new_Sorter100|16930_ ,
    \new_Sorter100|16931_ , \new_Sorter100|16932_ , \new_Sorter100|16933_ ,
    \new_Sorter100|16934_ , \new_Sorter100|16935_ , \new_Sorter100|16936_ ,
    \new_Sorter100|16937_ , \new_Sorter100|16938_ , \new_Sorter100|16939_ ,
    \new_Sorter100|16940_ , \new_Sorter100|16941_ , \new_Sorter100|16942_ ,
    \new_Sorter100|16943_ , \new_Sorter100|16944_ , \new_Sorter100|16945_ ,
    \new_Sorter100|16946_ , \new_Sorter100|16947_ , \new_Sorter100|16948_ ,
    \new_Sorter100|16949_ , \new_Sorter100|16950_ , \new_Sorter100|16951_ ,
    \new_Sorter100|16952_ , \new_Sorter100|16953_ , \new_Sorter100|16954_ ,
    \new_Sorter100|16955_ , \new_Sorter100|16956_ , \new_Sorter100|16957_ ,
    \new_Sorter100|16958_ , \new_Sorter100|16959_ , \new_Sorter100|16960_ ,
    \new_Sorter100|16961_ , \new_Sorter100|16962_ , \new_Sorter100|16963_ ,
    \new_Sorter100|16964_ , \new_Sorter100|16965_ , \new_Sorter100|16966_ ,
    \new_Sorter100|16967_ , \new_Sorter100|16968_ , \new_Sorter100|16969_ ,
    \new_Sorter100|16970_ , \new_Sorter100|16971_ , \new_Sorter100|16972_ ,
    \new_Sorter100|16973_ , \new_Sorter100|16974_ , \new_Sorter100|16975_ ,
    \new_Sorter100|16976_ , \new_Sorter100|16977_ , \new_Sorter100|16978_ ,
    \new_Sorter100|16979_ , \new_Sorter100|16980_ , \new_Sorter100|16981_ ,
    \new_Sorter100|16982_ , \new_Sorter100|16983_ , \new_Sorter100|16984_ ,
    \new_Sorter100|16985_ , \new_Sorter100|16986_ , \new_Sorter100|16987_ ,
    \new_Sorter100|16988_ , \new_Sorter100|16989_ , \new_Sorter100|16990_ ,
    \new_Sorter100|16991_ , \new_Sorter100|16992_ , \new_Sorter100|16993_ ,
    \new_Sorter100|16994_ , \new_Sorter100|16995_ , \new_Sorter100|16996_ ,
    \new_Sorter100|16997_ , \new_Sorter100|16998_ , \new_Sorter100|17000_ ,
    \new_Sorter100|17001_ , \new_Sorter100|17002_ , \new_Sorter100|17003_ ,
    \new_Sorter100|17004_ , \new_Sorter100|17005_ , \new_Sorter100|17006_ ,
    \new_Sorter100|17007_ , \new_Sorter100|17008_ , \new_Sorter100|17009_ ,
    \new_Sorter100|17010_ , \new_Sorter100|17011_ , \new_Sorter100|17012_ ,
    \new_Sorter100|17013_ , \new_Sorter100|17014_ , \new_Sorter100|17015_ ,
    \new_Sorter100|17016_ , \new_Sorter100|17017_ , \new_Sorter100|17018_ ,
    \new_Sorter100|17019_ , \new_Sorter100|17020_ , \new_Sorter100|17021_ ,
    \new_Sorter100|17022_ , \new_Sorter100|17023_ , \new_Sorter100|17024_ ,
    \new_Sorter100|17025_ , \new_Sorter100|17026_ , \new_Sorter100|17027_ ,
    \new_Sorter100|17028_ , \new_Sorter100|17029_ , \new_Sorter100|17030_ ,
    \new_Sorter100|17031_ , \new_Sorter100|17032_ , \new_Sorter100|17033_ ,
    \new_Sorter100|17034_ , \new_Sorter100|17035_ , \new_Sorter100|17036_ ,
    \new_Sorter100|17037_ , \new_Sorter100|17038_ , \new_Sorter100|17039_ ,
    \new_Sorter100|17040_ , \new_Sorter100|17041_ , \new_Sorter100|17042_ ,
    \new_Sorter100|17043_ , \new_Sorter100|17044_ , \new_Sorter100|17045_ ,
    \new_Sorter100|17046_ , \new_Sorter100|17047_ , \new_Sorter100|17048_ ,
    \new_Sorter100|17049_ , \new_Sorter100|17050_ , \new_Sorter100|17051_ ,
    \new_Sorter100|17052_ , \new_Sorter100|17053_ , \new_Sorter100|17054_ ,
    \new_Sorter100|17055_ , \new_Sorter100|17056_ , \new_Sorter100|17057_ ,
    \new_Sorter100|17058_ , \new_Sorter100|17059_ , \new_Sorter100|17060_ ,
    \new_Sorter100|17061_ , \new_Sorter100|17062_ , \new_Sorter100|17063_ ,
    \new_Sorter100|17064_ , \new_Sorter100|17065_ , \new_Sorter100|17066_ ,
    \new_Sorter100|17067_ , \new_Sorter100|17068_ , \new_Sorter100|17069_ ,
    \new_Sorter100|17070_ , \new_Sorter100|17071_ , \new_Sorter100|17072_ ,
    \new_Sorter100|17073_ , \new_Sorter100|17074_ , \new_Sorter100|17075_ ,
    \new_Sorter100|17076_ , \new_Sorter100|17077_ , \new_Sorter100|17078_ ,
    \new_Sorter100|17079_ , \new_Sorter100|17080_ , \new_Sorter100|17081_ ,
    \new_Sorter100|17082_ , \new_Sorter100|17083_ , \new_Sorter100|17084_ ,
    \new_Sorter100|17085_ , \new_Sorter100|17086_ , \new_Sorter100|17087_ ,
    \new_Sorter100|17088_ , \new_Sorter100|17089_ , \new_Sorter100|17090_ ,
    \new_Sorter100|17091_ , \new_Sorter100|17092_ , \new_Sorter100|17093_ ,
    \new_Sorter100|17094_ , \new_Sorter100|17095_ , \new_Sorter100|17096_ ,
    \new_Sorter100|17097_ , \new_Sorter100|17098_ , \new_Sorter100|17099_ ,
    \new_Sorter100|17100_ , \new_Sorter100|17199_ , \new_Sorter100|17101_ ,
    \new_Sorter100|17102_ , \new_Sorter100|17103_ , \new_Sorter100|17104_ ,
    \new_Sorter100|17105_ , \new_Sorter100|17106_ , \new_Sorter100|17107_ ,
    \new_Sorter100|17108_ , \new_Sorter100|17109_ , \new_Sorter100|17110_ ,
    \new_Sorter100|17111_ , \new_Sorter100|17112_ , \new_Sorter100|17113_ ,
    \new_Sorter100|17114_ , \new_Sorter100|17115_ , \new_Sorter100|17116_ ,
    \new_Sorter100|17117_ , \new_Sorter100|17118_ , \new_Sorter100|17119_ ,
    \new_Sorter100|17120_ , \new_Sorter100|17121_ , \new_Sorter100|17122_ ,
    \new_Sorter100|17123_ , \new_Sorter100|17124_ , \new_Sorter100|17125_ ,
    \new_Sorter100|17126_ , \new_Sorter100|17127_ , \new_Sorter100|17128_ ,
    \new_Sorter100|17129_ , \new_Sorter100|17130_ , \new_Sorter100|17131_ ,
    \new_Sorter100|17132_ , \new_Sorter100|17133_ , \new_Sorter100|17134_ ,
    \new_Sorter100|17135_ , \new_Sorter100|17136_ , \new_Sorter100|17137_ ,
    \new_Sorter100|17138_ , \new_Sorter100|17139_ , \new_Sorter100|17140_ ,
    \new_Sorter100|17141_ , \new_Sorter100|17142_ , \new_Sorter100|17143_ ,
    \new_Sorter100|17144_ , \new_Sorter100|17145_ , \new_Sorter100|17146_ ,
    \new_Sorter100|17147_ , \new_Sorter100|17148_ , \new_Sorter100|17149_ ,
    \new_Sorter100|17150_ , \new_Sorter100|17151_ , \new_Sorter100|17152_ ,
    \new_Sorter100|17153_ , \new_Sorter100|17154_ , \new_Sorter100|17155_ ,
    \new_Sorter100|17156_ , \new_Sorter100|17157_ , \new_Sorter100|17158_ ,
    \new_Sorter100|17159_ , \new_Sorter100|17160_ , \new_Sorter100|17161_ ,
    \new_Sorter100|17162_ , \new_Sorter100|17163_ , \new_Sorter100|17164_ ,
    \new_Sorter100|17165_ , \new_Sorter100|17166_ , \new_Sorter100|17167_ ,
    \new_Sorter100|17168_ , \new_Sorter100|17169_ , \new_Sorter100|17170_ ,
    \new_Sorter100|17171_ , \new_Sorter100|17172_ , \new_Sorter100|17173_ ,
    \new_Sorter100|17174_ , \new_Sorter100|17175_ , \new_Sorter100|17176_ ,
    \new_Sorter100|17177_ , \new_Sorter100|17178_ , \new_Sorter100|17179_ ,
    \new_Sorter100|17180_ , \new_Sorter100|17181_ , \new_Sorter100|17182_ ,
    \new_Sorter100|17183_ , \new_Sorter100|17184_ , \new_Sorter100|17185_ ,
    \new_Sorter100|17186_ , \new_Sorter100|17187_ , \new_Sorter100|17188_ ,
    \new_Sorter100|17189_ , \new_Sorter100|17190_ , \new_Sorter100|17191_ ,
    \new_Sorter100|17192_ , \new_Sorter100|17193_ , \new_Sorter100|17194_ ,
    \new_Sorter100|17195_ , \new_Sorter100|17196_ , \new_Sorter100|17197_ ,
    \new_Sorter100|17198_ , \new_Sorter100|17200_ , \new_Sorter100|17201_ ,
    \new_Sorter100|17202_ , \new_Sorter100|17203_ , \new_Sorter100|17204_ ,
    \new_Sorter100|17205_ , \new_Sorter100|17206_ , \new_Sorter100|17207_ ,
    \new_Sorter100|17208_ , \new_Sorter100|17209_ , \new_Sorter100|17210_ ,
    \new_Sorter100|17211_ , \new_Sorter100|17212_ , \new_Sorter100|17213_ ,
    \new_Sorter100|17214_ , \new_Sorter100|17215_ , \new_Sorter100|17216_ ,
    \new_Sorter100|17217_ , \new_Sorter100|17218_ , \new_Sorter100|17219_ ,
    \new_Sorter100|17220_ , \new_Sorter100|17221_ , \new_Sorter100|17222_ ,
    \new_Sorter100|17223_ , \new_Sorter100|17224_ , \new_Sorter100|17225_ ,
    \new_Sorter100|17226_ , \new_Sorter100|17227_ , \new_Sorter100|17228_ ,
    \new_Sorter100|17229_ , \new_Sorter100|17230_ , \new_Sorter100|17231_ ,
    \new_Sorter100|17232_ , \new_Sorter100|17233_ , \new_Sorter100|17234_ ,
    \new_Sorter100|17235_ , \new_Sorter100|17236_ , \new_Sorter100|17237_ ,
    \new_Sorter100|17238_ , \new_Sorter100|17239_ , \new_Sorter100|17240_ ,
    \new_Sorter100|17241_ , \new_Sorter100|17242_ , \new_Sorter100|17243_ ,
    \new_Sorter100|17244_ , \new_Sorter100|17245_ , \new_Sorter100|17246_ ,
    \new_Sorter100|17247_ , \new_Sorter100|17248_ , \new_Sorter100|17249_ ,
    \new_Sorter100|17250_ , \new_Sorter100|17251_ , \new_Sorter100|17252_ ,
    \new_Sorter100|17253_ , \new_Sorter100|17254_ , \new_Sorter100|17255_ ,
    \new_Sorter100|17256_ , \new_Sorter100|17257_ , \new_Sorter100|17258_ ,
    \new_Sorter100|17259_ , \new_Sorter100|17260_ , \new_Sorter100|17261_ ,
    \new_Sorter100|17262_ , \new_Sorter100|17263_ , \new_Sorter100|17264_ ,
    \new_Sorter100|17265_ , \new_Sorter100|17266_ , \new_Sorter100|17267_ ,
    \new_Sorter100|17268_ , \new_Sorter100|17269_ , \new_Sorter100|17270_ ,
    \new_Sorter100|17271_ , \new_Sorter100|17272_ , \new_Sorter100|17273_ ,
    \new_Sorter100|17274_ , \new_Sorter100|17275_ , \new_Sorter100|17276_ ,
    \new_Sorter100|17277_ , \new_Sorter100|17278_ , \new_Sorter100|17279_ ,
    \new_Sorter100|17280_ , \new_Sorter100|17281_ , \new_Sorter100|17282_ ,
    \new_Sorter100|17283_ , \new_Sorter100|17284_ , \new_Sorter100|17285_ ,
    \new_Sorter100|17286_ , \new_Sorter100|17287_ , \new_Sorter100|17288_ ,
    \new_Sorter100|17289_ , \new_Sorter100|17290_ , \new_Sorter100|17291_ ,
    \new_Sorter100|17292_ , \new_Sorter100|17293_ , \new_Sorter100|17294_ ,
    \new_Sorter100|17295_ , \new_Sorter100|17296_ , \new_Sorter100|17297_ ,
    \new_Sorter100|17298_ , \new_Sorter100|17299_ , \new_Sorter100|17300_ ,
    \new_Sorter100|17399_ , \new_Sorter100|17301_ , \new_Sorter100|17302_ ,
    \new_Sorter100|17303_ , \new_Sorter100|17304_ , \new_Sorter100|17305_ ,
    \new_Sorter100|17306_ , \new_Sorter100|17307_ , \new_Sorter100|17308_ ,
    \new_Sorter100|17309_ , \new_Sorter100|17310_ , \new_Sorter100|17311_ ,
    \new_Sorter100|17312_ , \new_Sorter100|17313_ , \new_Sorter100|17314_ ,
    \new_Sorter100|17315_ , \new_Sorter100|17316_ , \new_Sorter100|17317_ ,
    \new_Sorter100|17318_ , \new_Sorter100|17319_ , \new_Sorter100|17320_ ,
    \new_Sorter100|17321_ , \new_Sorter100|17322_ , \new_Sorter100|17323_ ,
    \new_Sorter100|17324_ , \new_Sorter100|17325_ , \new_Sorter100|17326_ ,
    \new_Sorter100|17327_ , \new_Sorter100|17328_ , \new_Sorter100|17329_ ,
    \new_Sorter100|17330_ , \new_Sorter100|17331_ , \new_Sorter100|17332_ ,
    \new_Sorter100|17333_ , \new_Sorter100|17334_ , \new_Sorter100|17335_ ,
    \new_Sorter100|17336_ , \new_Sorter100|17337_ , \new_Sorter100|17338_ ,
    \new_Sorter100|17339_ , \new_Sorter100|17340_ , \new_Sorter100|17341_ ,
    \new_Sorter100|17342_ , \new_Sorter100|17343_ , \new_Sorter100|17344_ ,
    \new_Sorter100|17345_ , \new_Sorter100|17346_ , \new_Sorter100|17347_ ,
    \new_Sorter100|17348_ , \new_Sorter100|17349_ , \new_Sorter100|17350_ ,
    \new_Sorter100|17351_ , \new_Sorter100|17352_ , \new_Sorter100|17353_ ,
    \new_Sorter100|17354_ , \new_Sorter100|17355_ , \new_Sorter100|17356_ ,
    \new_Sorter100|17357_ , \new_Sorter100|17358_ , \new_Sorter100|17359_ ,
    \new_Sorter100|17360_ , \new_Sorter100|17361_ , \new_Sorter100|17362_ ,
    \new_Sorter100|17363_ , \new_Sorter100|17364_ , \new_Sorter100|17365_ ,
    \new_Sorter100|17366_ , \new_Sorter100|17367_ , \new_Sorter100|17368_ ,
    \new_Sorter100|17369_ , \new_Sorter100|17370_ , \new_Sorter100|17371_ ,
    \new_Sorter100|17372_ , \new_Sorter100|17373_ , \new_Sorter100|17374_ ,
    \new_Sorter100|17375_ , \new_Sorter100|17376_ , \new_Sorter100|17377_ ,
    \new_Sorter100|17378_ , \new_Sorter100|17379_ , \new_Sorter100|17380_ ,
    \new_Sorter100|17381_ , \new_Sorter100|17382_ , \new_Sorter100|17383_ ,
    \new_Sorter100|17384_ , \new_Sorter100|17385_ , \new_Sorter100|17386_ ,
    \new_Sorter100|17387_ , \new_Sorter100|17388_ , \new_Sorter100|17389_ ,
    \new_Sorter100|17390_ , \new_Sorter100|17391_ , \new_Sorter100|17392_ ,
    \new_Sorter100|17393_ , \new_Sorter100|17394_ , \new_Sorter100|17395_ ,
    \new_Sorter100|17396_ , \new_Sorter100|17397_ , \new_Sorter100|17398_ ,
    \new_Sorter100|17400_ , \new_Sorter100|17401_ , \new_Sorter100|17402_ ,
    \new_Sorter100|17403_ , \new_Sorter100|17404_ , \new_Sorter100|17405_ ,
    \new_Sorter100|17406_ , \new_Sorter100|17407_ , \new_Sorter100|17408_ ,
    \new_Sorter100|17409_ , \new_Sorter100|17410_ , \new_Sorter100|17411_ ,
    \new_Sorter100|17412_ , \new_Sorter100|17413_ , \new_Sorter100|17414_ ,
    \new_Sorter100|17415_ , \new_Sorter100|17416_ , \new_Sorter100|17417_ ,
    \new_Sorter100|17418_ , \new_Sorter100|17419_ , \new_Sorter100|17420_ ,
    \new_Sorter100|17421_ , \new_Sorter100|17422_ , \new_Sorter100|17423_ ,
    \new_Sorter100|17424_ , \new_Sorter100|17425_ , \new_Sorter100|17426_ ,
    \new_Sorter100|17427_ , \new_Sorter100|17428_ , \new_Sorter100|17429_ ,
    \new_Sorter100|17430_ , \new_Sorter100|17431_ , \new_Sorter100|17432_ ,
    \new_Sorter100|17433_ , \new_Sorter100|17434_ , \new_Sorter100|17435_ ,
    \new_Sorter100|17436_ , \new_Sorter100|17437_ , \new_Sorter100|17438_ ,
    \new_Sorter100|17439_ , \new_Sorter100|17440_ , \new_Sorter100|17441_ ,
    \new_Sorter100|17442_ , \new_Sorter100|17443_ , \new_Sorter100|17444_ ,
    \new_Sorter100|17445_ , \new_Sorter100|17446_ , \new_Sorter100|17447_ ,
    \new_Sorter100|17448_ , \new_Sorter100|17449_ , \new_Sorter100|17450_ ,
    \new_Sorter100|17451_ , \new_Sorter100|17452_ , \new_Sorter100|17453_ ,
    \new_Sorter100|17454_ , \new_Sorter100|17455_ , \new_Sorter100|17456_ ,
    \new_Sorter100|17457_ , \new_Sorter100|17458_ , \new_Sorter100|17459_ ,
    \new_Sorter100|17460_ , \new_Sorter100|17461_ , \new_Sorter100|17462_ ,
    \new_Sorter100|17463_ , \new_Sorter100|17464_ , \new_Sorter100|17465_ ,
    \new_Sorter100|17466_ , \new_Sorter100|17467_ , \new_Sorter100|17468_ ,
    \new_Sorter100|17469_ , \new_Sorter100|17470_ , \new_Sorter100|17471_ ,
    \new_Sorter100|17472_ , \new_Sorter100|17473_ , \new_Sorter100|17474_ ,
    \new_Sorter100|17475_ , \new_Sorter100|17476_ , \new_Sorter100|17477_ ,
    \new_Sorter100|17478_ , \new_Sorter100|17479_ , \new_Sorter100|17480_ ,
    \new_Sorter100|17481_ , \new_Sorter100|17482_ , \new_Sorter100|17483_ ,
    \new_Sorter100|17484_ , \new_Sorter100|17485_ , \new_Sorter100|17486_ ,
    \new_Sorter100|17487_ , \new_Sorter100|17488_ , \new_Sorter100|17489_ ,
    \new_Sorter100|17490_ , \new_Sorter100|17491_ , \new_Sorter100|17492_ ,
    \new_Sorter100|17493_ , \new_Sorter100|17494_ , \new_Sorter100|17495_ ,
    \new_Sorter100|17496_ , \new_Sorter100|17497_ , \new_Sorter100|17498_ ,
    \new_Sorter100|17499_ , \new_Sorter100|17500_ , \new_Sorter100|17599_ ,
    \new_Sorter100|17501_ , \new_Sorter100|17502_ , \new_Sorter100|17503_ ,
    \new_Sorter100|17504_ , \new_Sorter100|17505_ , \new_Sorter100|17506_ ,
    \new_Sorter100|17507_ , \new_Sorter100|17508_ , \new_Sorter100|17509_ ,
    \new_Sorter100|17510_ , \new_Sorter100|17511_ , \new_Sorter100|17512_ ,
    \new_Sorter100|17513_ , \new_Sorter100|17514_ , \new_Sorter100|17515_ ,
    \new_Sorter100|17516_ , \new_Sorter100|17517_ , \new_Sorter100|17518_ ,
    \new_Sorter100|17519_ , \new_Sorter100|17520_ , \new_Sorter100|17521_ ,
    \new_Sorter100|17522_ , \new_Sorter100|17523_ , \new_Sorter100|17524_ ,
    \new_Sorter100|17525_ , \new_Sorter100|17526_ , \new_Sorter100|17527_ ,
    \new_Sorter100|17528_ , \new_Sorter100|17529_ , \new_Sorter100|17530_ ,
    \new_Sorter100|17531_ , \new_Sorter100|17532_ , \new_Sorter100|17533_ ,
    \new_Sorter100|17534_ , \new_Sorter100|17535_ , \new_Sorter100|17536_ ,
    \new_Sorter100|17537_ , \new_Sorter100|17538_ , \new_Sorter100|17539_ ,
    \new_Sorter100|17540_ , \new_Sorter100|17541_ , \new_Sorter100|17542_ ,
    \new_Sorter100|17543_ , \new_Sorter100|17544_ , \new_Sorter100|17545_ ,
    \new_Sorter100|17546_ , \new_Sorter100|17547_ , \new_Sorter100|17548_ ,
    \new_Sorter100|17549_ , \new_Sorter100|17550_ , \new_Sorter100|17551_ ,
    \new_Sorter100|17552_ , \new_Sorter100|17553_ , \new_Sorter100|17554_ ,
    \new_Sorter100|17555_ , \new_Sorter100|17556_ , \new_Sorter100|17557_ ,
    \new_Sorter100|17558_ , \new_Sorter100|17559_ , \new_Sorter100|17560_ ,
    \new_Sorter100|17561_ , \new_Sorter100|17562_ , \new_Sorter100|17563_ ,
    \new_Sorter100|17564_ , \new_Sorter100|17565_ , \new_Sorter100|17566_ ,
    \new_Sorter100|17567_ , \new_Sorter100|17568_ , \new_Sorter100|17569_ ,
    \new_Sorter100|17570_ , \new_Sorter100|17571_ , \new_Sorter100|17572_ ,
    \new_Sorter100|17573_ , \new_Sorter100|17574_ , \new_Sorter100|17575_ ,
    \new_Sorter100|17576_ , \new_Sorter100|17577_ , \new_Sorter100|17578_ ,
    \new_Sorter100|17579_ , \new_Sorter100|17580_ , \new_Sorter100|17581_ ,
    \new_Sorter100|17582_ , \new_Sorter100|17583_ , \new_Sorter100|17584_ ,
    \new_Sorter100|17585_ , \new_Sorter100|17586_ , \new_Sorter100|17587_ ,
    \new_Sorter100|17588_ , \new_Sorter100|17589_ , \new_Sorter100|17590_ ,
    \new_Sorter100|17591_ , \new_Sorter100|17592_ , \new_Sorter100|17593_ ,
    \new_Sorter100|17594_ , \new_Sorter100|17595_ , \new_Sorter100|17596_ ,
    \new_Sorter100|17597_ , \new_Sorter100|17598_ , \new_Sorter100|17600_ ,
    \new_Sorter100|17601_ , \new_Sorter100|17602_ , \new_Sorter100|17603_ ,
    \new_Sorter100|17604_ , \new_Sorter100|17605_ , \new_Sorter100|17606_ ,
    \new_Sorter100|17607_ , \new_Sorter100|17608_ , \new_Sorter100|17609_ ,
    \new_Sorter100|17610_ , \new_Sorter100|17611_ , \new_Sorter100|17612_ ,
    \new_Sorter100|17613_ , \new_Sorter100|17614_ , \new_Sorter100|17615_ ,
    \new_Sorter100|17616_ , \new_Sorter100|17617_ , \new_Sorter100|17618_ ,
    \new_Sorter100|17619_ , \new_Sorter100|17620_ , \new_Sorter100|17621_ ,
    \new_Sorter100|17622_ , \new_Sorter100|17623_ , \new_Sorter100|17624_ ,
    \new_Sorter100|17625_ , \new_Sorter100|17626_ , \new_Sorter100|17627_ ,
    \new_Sorter100|17628_ , \new_Sorter100|17629_ , \new_Sorter100|17630_ ,
    \new_Sorter100|17631_ , \new_Sorter100|17632_ , \new_Sorter100|17633_ ,
    \new_Sorter100|17634_ , \new_Sorter100|17635_ , \new_Sorter100|17636_ ,
    \new_Sorter100|17637_ , \new_Sorter100|17638_ , \new_Sorter100|17639_ ,
    \new_Sorter100|17640_ , \new_Sorter100|17641_ , \new_Sorter100|17642_ ,
    \new_Sorter100|17643_ , \new_Sorter100|17644_ , \new_Sorter100|17645_ ,
    \new_Sorter100|17646_ , \new_Sorter100|17647_ , \new_Sorter100|17648_ ,
    \new_Sorter100|17649_ , \new_Sorter100|17650_ , \new_Sorter100|17651_ ,
    \new_Sorter100|17652_ , \new_Sorter100|17653_ , \new_Sorter100|17654_ ,
    \new_Sorter100|17655_ , \new_Sorter100|17656_ , \new_Sorter100|17657_ ,
    \new_Sorter100|17658_ , \new_Sorter100|17659_ , \new_Sorter100|17660_ ,
    \new_Sorter100|17661_ , \new_Sorter100|17662_ , \new_Sorter100|17663_ ,
    \new_Sorter100|17664_ , \new_Sorter100|17665_ , \new_Sorter100|17666_ ,
    \new_Sorter100|17667_ , \new_Sorter100|17668_ , \new_Sorter100|17669_ ,
    \new_Sorter100|17670_ , \new_Sorter100|17671_ , \new_Sorter100|17672_ ,
    \new_Sorter100|17673_ , \new_Sorter100|17674_ , \new_Sorter100|17675_ ,
    \new_Sorter100|17676_ , \new_Sorter100|17677_ , \new_Sorter100|17678_ ,
    \new_Sorter100|17679_ , \new_Sorter100|17680_ , \new_Sorter100|17681_ ,
    \new_Sorter100|17682_ , \new_Sorter100|17683_ , \new_Sorter100|17684_ ,
    \new_Sorter100|17685_ , \new_Sorter100|17686_ , \new_Sorter100|17687_ ,
    \new_Sorter100|17688_ , \new_Sorter100|17689_ , \new_Sorter100|17690_ ,
    \new_Sorter100|17691_ , \new_Sorter100|17692_ , \new_Sorter100|17693_ ,
    \new_Sorter100|17694_ , \new_Sorter100|17695_ , \new_Sorter100|17696_ ,
    \new_Sorter100|17697_ , \new_Sorter100|17698_ , \new_Sorter100|17699_ ,
    \new_Sorter100|17700_ , \new_Sorter100|17799_ , \new_Sorter100|17701_ ,
    \new_Sorter100|17702_ , \new_Sorter100|17703_ , \new_Sorter100|17704_ ,
    \new_Sorter100|17705_ , \new_Sorter100|17706_ , \new_Sorter100|17707_ ,
    \new_Sorter100|17708_ , \new_Sorter100|17709_ , \new_Sorter100|17710_ ,
    \new_Sorter100|17711_ , \new_Sorter100|17712_ , \new_Sorter100|17713_ ,
    \new_Sorter100|17714_ , \new_Sorter100|17715_ , \new_Sorter100|17716_ ,
    \new_Sorter100|17717_ , \new_Sorter100|17718_ , \new_Sorter100|17719_ ,
    \new_Sorter100|17720_ , \new_Sorter100|17721_ , \new_Sorter100|17722_ ,
    \new_Sorter100|17723_ , \new_Sorter100|17724_ , \new_Sorter100|17725_ ,
    \new_Sorter100|17726_ , \new_Sorter100|17727_ , \new_Sorter100|17728_ ,
    \new_Sorter100|17729_ , \new_Sorter100|17730_ , \new_Sorter100|17731_ ,
    \new_Sorter100|17732_ , \new_Sorter100|17733_ , \new_Sorter100|17734_ ,
    \new_Sorter100|17735_ , \new_Sorter100|17736_ , \new_Sorter100|17737_ ,
    \new_Sorter100|17738_ , \new_Sorter100|17739_ , \new_Sorter100|17740_ ,
    \new_Sorter100|17741_ , \new_Sorter100|17742_ , \new_Sorter100|17743_ ,
    \new_Sorter100|17744_ , \new_Sorter100|17745_ , \new_Sorter100|17746_ ,
    \new_Sorter100|17747_ , \new_Sorter100|17748_ , \new_Sorter100|17749_ ,
    \new_Sorter100|17750_ , \new_Sorter100|17751_ , \new_Sorter100|17752_ ,
    \new_Sorter100|17753_ , \new_Sorter100|17754_ , \new_Sorter100|17755_ ,
    \new_Sorter100|17756_ , \new_Sorter100|17757_ , \new_Sorter100|17758_ ,
    \new_Sorter100|17759_ , \new_Sorter100|17760_ , \new_Sorter100|17761_ ,
    \new_Sorter100|17762_ , \new_Sorter100|17763_ , \new_Sorter100|17764_ ,
    \new_Sorter100|17765_ , \new_Sorter100|17766_ , \new_Sorter100|17767_ ,
    \new_Sorter100|17768_ , \new_Sorter100|17769_ , \new_Sorter100|17770_ ,
    \new_Sorter100|17771_ , \new_Sorter100|17772_ , \new_Sorter100|17773_ ,
    \new_Sorter100|17774_ , \new_Sorter100|17775_ , \new_Sorter100|17776_ ,
    \new_Sorter100|17777_ , \new_Sorter100|17778_ , \new_Sorter100|17779_ ,
    \new_Sorter100|17780_ , \new_Sorter100|17781_ , \new_Sorter100|17782_ ,
    \new_Sorter100|17783_ , \new_Sorter100|17784_ , \new_Sorter100|17785_ ,
    \new_Sorter100|17786_ , \new_Sorter100|17787_ , \new_Sorter100|17788_ ,
    \new_Sorter100|17789_ , \new_Sorter100|17790_ , \new_Sorter100|17791_ ,
    \new_Sorter100|17792_ , \new_Sorter100|17793_ , \new_Sorter100|17794_ ,
    \new_Sorter100|17795_ , \new_Sorter100|17796_ , \new_Sorter100|17797_ ,
    \new_Sorter100|17798_ , \new_Sorter100|17800_ , \new_Sorter100|17801_ ,
    \new_Sorter100|17802_ , \new_Sorter100|17803_ , \new_Sorter100|17804_ ,
    \new_Sorter100|17805_ , \new_Sorter100|17806_ , \new_Sorter100|17807_ ,
    \new_Sorter100|17808_ , \new_Sorter100|17809_ , \new_Sorter100|17810_ ,
    \new_Sorter100|17811_ , \new_Sorter100|17812_ , \new_Sorter100|17813_ ,
    \new_Sorter100|17814_ , \new_Sorter100|17815_ , \new_Sorter100|17816_ ,
    \new_Sorter100|17817_ , \new_Sorter100|17818_ , \new_Sorter100|17819_ ,
    \new_Sorter100|17820_ , \new_Sorter100|17821_ , \new_Sorter100|17822_ ,
    \new_Sorter100|17823_ , \new_Sorter100|17824_ , \new_Sorter100|17825_ ,
    \new_Sorter100|17826_ , \new_Sorter100|17827_ , \new_Sorter100|17828_ ,
    \new_Sorter100|17829_ , \new_Sorter100|17830_ , \new_Sorter100|17831_ ,
    \new_Sorter100|17832_ , \new_Sorter100|17833_ , \new_Sorter100|17834_ ,
    \new_Sorter100|17835_ , \new_Sorter100|17836_ , \new_Sorter100|17837_ ,
    \new_Sorter100|17838_ , \new_Sorter100|17839_ , \new_Sorter100|17840_ ,
    \new_Sorter100|17841_ , \new_Sorter100|17842_ , \new_Sorter100|17843_ ,
    \new_Sorter100|17844_ , \new_Sorter100|17845_ , \new_Sorter100|17846_ ,
    \new_Sorter100|17847_ , \new_Sorter100|17848_ , \new_Sorter100|17849_ ,
    \new_Sorter100|17850_ , \new_Sorter100|17851_ , \new_Sorter100|17852_ ,
    \new_Sorter100|17853_ , \new_Sorter100|17854_ , \new_Sorter100|17855_ ,
    \new_Sorter100|17856_ , \new_Sorter100|17857_ , \new_Sorter100|17858_ ,
    \new_Sorter100|17859_ , \new_Sorter100|17860_ , \new_Sorter100|17861_ ,
    \new_Sorter100|17862_ , \new_Sorter100|17863_ , \new_Sorter100|17864_ ,
    \new_Sorter100|17865_ , \new_Sorter100|17866_ , \new_Sorter100|17867_ ,
    \new_Sorter100|17868_ , \new_Sorter100|17869_ , \new_Sorter100|17870_ ,
    \new_Sorter100|17871_ , \new_Sorter100|17872_ , \new_Sorter100|17873_ ,
    \new_Sorter100|17874_ , \new_Sorter100|17875_ , \new_Sorter100|17876_ ,
    \new_Sorter100|17877_ , \new_Sorter100|17878_ , \new_Sorter100|17879_ ,
    \new_Sorter100|17880_ , \new_Sorter100|17881_ , \new_Sorter100|17882_ ,
    \new_Sorter100|17883_ , \new_Sorter100|17884_ , \new_Sorter100|17885_ ,
    \new_Sorter100|17886_ , \new_Sorter100|17887_ , \new_Sorter100|17888_ ,
    \new_Sorter100|17889_ , \new_Sorter100|17890_ , \new_Sorter100|17891_ ,
    \new_Sorter100|17892_ , \new_Sorter100|17893_ , \new_Sorter100|17894_ ,
    \new_Sorter100|17895_ , \new_Sorter100|17896_ , \new_Sorter100|17897_ ,
    \new_Sorter100|17898_ , \new_Sorter100|17899_ , \new_Sorter100|17900_ ,
    \new_Sorter100|17999_ , \new_Sorter100|17901_ , \new_Sorter100|17902_ ,
    \new_Sorter100|17903_ , \new_Sorter100|17904_ , \new_Sorter100|17905_ ,
    \new_Sorter100|17906_ , \new_Sorter100|17907_ , \new_Sorter100|17908_ ,
    \new_Sorter100|17909_ , \new_Sorter100|17910_ , \new_Sorter100|17911_ ,
    \new_Sorter100|17912_ , \new_Sorter100|17913_ , \new_Sorter100|17914_ ,
    \new_Sorter100|17915_ , \new_Sorter100|17916_ , \new_Sorter100|17917_ ,
    \new_Sorter100|17918_ , \new_Sorter100|17919_ , \new_Sorter100|17920_ ,
    \new_Sorter100|17921_ , \new_Sorter100|17922_ , \new_Sorter100|17923_ ,
    \new_Sorter100|17924_ , \new_Sorter100|17925_ , \new_Sorter100|17926_ ,
    \new_Sorter100|17927_ , \new_Sorter100|17928_ , \new_Sorter100|17929_ ,
    \new_Sorter100|17930_ , \new_Sorter100|17931_ , \new_Sorter100|17932_ ,
    \new_Sorter100|17933_ , \new_Sorter100|17934_ , \new_Sorter100|17935_ ,
    \new_Sorter100|17936_ , \new_Sorter100|17937_ , \new_Sorter100|17938_ ,
    \new_Sorter100|17939_ , \new_Sorter100|17940_ , \new_Sorter100|17941_ ,
    \new_Sorter100|17942_ , \new_Sorter100|17943_ , \new_Sorter100|17944_ ,
    \new_Sorter100|17945_ , \new_Sorter100|17946_ , \new_Sorter100|17947_ ,
    \new_Sorter100|17948_ , \new_Sorter100|17949_ , \new_Sorter100|17950_ ,
    \new_Sorter100|17951_ , \new_Sorter100|17952_ , \new_Sorter100|17953_ ,
    \new_Sorter100|17954_ , \new_Sorter100|17955_ , \new_Sorter100|17956_ ,
    \new_Sorter100|17957_ , \new_Sorter100|17958_ , \new_Sorter100|17959_ ,
    \new_Sorter100|17960_ , \new_Sorter100|17961_ , \new_Sorter100|17962_ ,
    \new_Sorter100|17963_ , \new_Sorter100|17964_ , \new_Sorter100|17965_ ,
    \new_Sorter100|17966_ , \new_Sorter100|17967_ , \new_Sorter100|17968_ ,
    \new_Sorter100|17969_ , \new_Sorter100|17970_ , \new_Sorter100|17971_ ,
    \new_Sorter100|17972_ , \new_Sorter100|17973_ , \new_Sorter100|17974_ ,
    \new_Sorter100|17975_ , \new_Sorter100|17976_ , \new_Sorter100|17977_ ,
    \new_Sorter100|17978_ , \new_Sorter100|17979_ , \new_Sorter100|17980_ ,
    \new_Sorter100|17981_ , \new_Sorter100|17982_ , \new_Sorter100|17983_ ,
    \new_Sorter100|17984_ , \new_Sorter100|17985_ , \new_Sorter100|17986_ ,
    \new_Sorter100|17987_ , \new_Sorter100|17988_ , \new_Sorter100|17989_ ,
    \new_Sorter100|17990_ , \new_Sorter100|17991_ , \new_Sorter100|17992_ ,
    \new_Sorter100|17993_ , \new_Sorter100|17994_ , \new_Sorter100|17995_ ,
    \new_Sorter100|17996_ , \new_Sorter100|17997_ , \new_Sorter100|17998_ ,
    \new_Sorter100|18000_ , \new_Sorter100|18001_ , \new_Sorter100|18002_ ,
    \new_Sorter100|18003_ , \new_Sorter100|18004_ , \new_Sorter100|18005_ ,
    \new_Sorter100|18006_ , \new_Sorter100|18007_ , \new_Sorter100|18008_ ,
    \new_Sorter100|18009_ , \new_Sorter100|18010_ , \new_Sorter100|18011_ ,
    \new_Sorter100|18012_ , \new_Sorter100|18013_ , \new_Sorter100|18014_ ,
    \new_Sorter100|18015_ , \new_Sorter100|18016_ , \new_Sorter100|18017_ ,
    \new_Sorter100|18018_ , \new_Sorter100|18019_ , \new_Sorter100|18020_ ,
    \new_Sorter100|18021_ , \new_Sorter100|18022_ , \new_Sorter100|18023_ ,
    \new_Sorter100|18024_ , \new_Sorter100|18025_ , \new_Sorter100|18026_ ,
    \new_Sorter100|18027_ , \new_Sorter100|18028_ , \new_Sorter100|18029_ ,
    \new_Sorter100|18030_ , \new_Sorter100|18031_ , \new_Sorter100|18032_ ,
    \new_Sorter100|18033_ , \new_Sorter100|18034_ , \new_Sorter100|18035_ ,
    \new_Sorter100|18036_ , \new_Sorter100|18037_ , \new_Sorter100|18038_ ,
    \new_Sorter100|18039_ , \new_Sorter100|18040_ , \new_Sorter100|18041_ ,
    \new_Sorter100|18042_ , \new_Sorter100|18043_ , \new_Sorter100|18044_ ,
    \new_Sorter100|18045_ , \new_Sorter100|18046_ , \new_Sorter100|18047_ ,
    \new_Sorter100|18048_ , \new_Sorter100|18049_ , \new_Sorter100|18050_ ,
    \new_Sorter100|18051_ , \new_Sorter100|18052_ , \new_Sorter100|18053_ ,
    \new_Sorter100|18054_ , \new_Sorter100|18055_ , \new_Sorter100|18056_ ,
    \new_Sorter100|18057_ , \new_Sorter100|18058_ , \new_Sorter100|18059_ ,
    \new_Sorter100|18060_ , \new_Sorter100|18061_ , \new_Sorter100|18062_ ,
    \new_Sorter100|18063_ , \new_Sorter100|18064_ , \new_Sorter100|18065_ ,
    \new_Sorter100|18066_ , \new_Sorter100|18067_ , \new_Sorter100|18068_ ,
    \new_Sorter100|18069_ , \new_Sorter100|18070_ , \new_Sorter100|18071_ ,
    \new_Sorter100|18072_ , \new_Sorter100|18073_ , \new_Sorter100|18074_ ,
    \new_Sorter100|18075_ , \new_Sorter100|18076_ , \new_Sorter100|18077_ ,
    \new_Sorter100|18078_ , \new_Sorter100|18079_ , \new_Sorter100|18080_ ,
    \new_Sorter100|18081_ , \new_Sorter100|18082_ , \new_Sorter100|18083_ ,
    \new_Sorter100|18084_ , \new_Sorter100|18085_ , \new_Sorter100|18086_ ,
    \new_Sorter100|18087_ , \new_Sorter100|18088_ , \new_Sorter100|18089_ ,
    \new_Sorter100|18090_ , \new_Sorter100|18091_ , \new_Sorter100|18092_ ,
    \new_Sorter100|18093_ , \new_Sorter100|18094_ , \new_Sorter100|18095_ ,
    \new_Sorter100|18096_ , \new_Sorter100|18097_ , \new_Sorter100|18098_ ,
    \new_Sorter100|18099_ , \new_Sorter100|18100_ , \new_Sorter100|18199_ ,
    \new_Sorter100|18101_ , \new_Sorter100|18102_ , \new_Sorter100|18103_ ,
    \new_Sorter100|18104_ , \new_Sorter100|18105_ , \new_Sorter100|18106_ ,
    \new_Sorter100|18107_ , \new_Sorter100|18108_ , \new_Sorter100|18109_ ,
    \new_Sorter100|18110_ , \new_Sorter100|18111_ , \new_Sorter100|18112_ ,
    \new_Sorter100|18113_ , \new_Sorter100|18114_ , \new_Sorter100|18115_ ,
    \new_Sorter100|18116_ , \new_Sorter100|18117_ , \new_Sorter100|18118_ ,
    \new_Sorter100|18119_ , \new_Sorter100|18120_ , \new_Sorter100|18121_ ,
    \new_Sorter100|18122_ , \new_Sorter100|18123_ , \new_Sorter100|18124_ ,
    \new_Sorter100|18125_ , \new_Sorter100|18126_ , \new_Sorter100|18127_ ,
    \new_Sorter100|18128_ , \new_Sorter100|18129_ , \new_Sorter100|18130_ ,
    \new_Sorter100|18131_ , \new_Sorter100|18132_ , \new_Sorter100|18133_ ,
    \new_Sorter100|18134_ , \new_Sorter100|18135_ , \new_Sorter100|18136_ ,
    \new_Sorter100|18137_ , \new_Sorter100|18138_ , \new_Sorter100|18139_ ,
    \new_Sorter100|18140_ , \new_Sorter100|18141_ , \new_Sorter100|18142_ ,
    \new_Sorter100|18143_ , \new_Sorter100|18144_ , \new_Sorter100|18145_ ,
    \new_Sorter100|18146_ , \new_Sorter100|18147_ , \new_Sorter100|18148_ ,
    \new_Sorter100|18149_ , \new_Sorter100|18150_ , \new_Sorter100|18151_ ,
    \new_Sorter100|18152_ , \new_Sorter100|18153_ , \new_Sorter100|18154_ ,
    \new_Sorter100|18155_ , \new_Sorter100|18156_ , \new_Sorter100|18157_ ,
    \new_Sorter100|18158_ , \new_Sorter100|18159_ , \new_Sorter100|18160_ ,
    \new_Sorter100|18161_ , \new_Sorter100|18162_ , \new_Sorter100|18163_ ,
    \new_Sorter100|18164_ , \new_Sorter100|18165_ , \new_Sorter100|18166_ ,
    \new_Sorter100|18167_ , \new_Sorter100|18168_ , \new_Sorter100|18169_ ,
    \new_Sorter100|18170_ , \new_Sorter100|18171_ , \new_Sorter100|18172_ ,
    \new_Sorter100|18173_ , \new_Sorter100|18174_ , \new_Sorter100|18175_ ,
    \new_Sorter100|18176_ , \new_Sorter100|18177_ , \new_Sorter100|18178_ ,
    \new_Sorter100|18179_ , \new_Sorter100|18180_ , \new_Sorter100|18181_ ,
    \new_Sorter100|18182_ , \new_Sorter100|18183_ , \new_Sorter100|18184_ ,
    \new_Sorter100|18185_ , \new_Sorter100|18186_ , \new_Sorter100|18187_ ,
    \new_Sorter100|18188_ , \new_Sorter100|18189_ , \new_Sorter100|18190_ ,
    \new_Sorter100|18191_ , \new_Sorter100|18192_ , \new_Sorter100|18193_ ,
    \new_Sorter100|18194_ , \new_Sorter100|18195_ , \new_Sorter100|18196_ ,
    \new_Sorter100|18197_ , \new_Sorter100|18198_ , \new_Sorter100|18200_ ,
    \new_Sorter100|18201_ , \new_Sorter100|18202_ , \new_Sorter100|18203_ ,
    \new_Sorter100|18204_ , \new_Sorter100|18205_ , \new_Sorter100|18206_ ,
    \new_Sorter100|18207_ , \new_Sorter100|18208_ , \new_Sorter100|18209_ ,
    \new_Sorter100|18210_ , \new_Sorter100|18211_ , \new_Sorter100|18212_ ,
    \new_Sorter100|18213_ , \new_Sorter100|18214_ , \new_Sorter100|18215_ ,
    \new_Sorter100|18216_ , \new_Sorter100|18217_ , \new_Sorter100|18218_ ,
    \new_Sorter100|18219_ , \new_Sorter100|18220_ , \new_Sorter100|18221_ ,
    \new_Sorter100|18222_ , \new_Sorter100|18223_ , \new_Sorter100|18224_ ,
    \new_Sorter100|18225_ , \new_Sorter100|18226_ , \new_Sorter100|18227_ ,
    \new_Sorter100|18228_ , \new_Sorter100|18229_ , \new_Sorter100|18230_ ,
    \new_Sorter100|18231_ , \new_Sorter100|18232_ , \new_Sorter100|18233_ ,
    \new_Sorter100|18234_ , \new_Sorter100|18235_ , \new_Sorter100|18236_ ,
    \new_Sorter100|18237_ , \new_Sorter100|18238_ , \new_Sorter100|18239_ ,
    \new_Sorter100|18240_ , \new_Sorter100|18241_ , \new_Sorter100|18242_ ,
    \new_Sorter100|18243_ , \new_Sorter100|18244_ , \new_Sorter100|18245_ ,
    \new_Sorter100|18246_ , \new_Sorter100|18247_ , \new_Sorter100|18248_ ,
    \new_Sorter100|18249_ , \new_Sorter100|18250_ , \new_Sorter100|18251_ ,
    \new_Sorter100|18252_ , \new_Sorter100|18253_ , \new_Sorter100|18254_ ,
    \new_Sorter100|18255_ , \new_Sorter100|18256_ , \new_Sorter100|18257_ ,
    \new_Sorter100|18258_ , \new_Sorter100|18259_ , \new_Sorter100|18260_ ,
    \new_Sorter100|18261_ , \new_Sorter100|18262_ , \new_Sorter100|18263_ ,
    \new_Sorter100|18264_ , \new_Sorter100|18265_ , \new_Sorter100|18266_ ,
    \new_Sorter100|18267_ , \new_Sorter100|18268_ , \new_Sorter100|18269_ ,
    \new_Sorter100|18270_ , \new_Sorter100|18271_ , \new_Sorter100|18272_ ,
    \new_Sorter100|18273_ , \new_Sorter100|18274_ , \new_Sorter100|18275_ ,
    \new_Sorter100|18276_ , \new_Sorter100|18277_ , \new_Sorter100|18278_ ,
    \new_Sorter100|18279_ , \new_Sorter100|18280_ , \new_Sorter100|18281_ ,
    \new_Sorter100|18282_ , \new_Sorter100|18283_ , \new_Sorter100|18284_ ,
    \new_Sorter100|18285_ , \new_Sorter100|18286_ , \new_Sorter100|18287_ ,
    \new_Sorter100|18288_ , \new_Sorter100|18289_ , \new_Sorter100|18290_ ,
    \new_Sorter100|18291_ , \new_Sorter100|18292_ , \new_Sorter100|18293_ ,
    \new_Sorter100|18294_ , \new_Sorter100|18295_ , \new_Sorter100|18296_ ,
    \new_Sorter100|18297_ , \new_Sorter100|18298_ , \new_Sorter100|18299_ ,
    \new_Sorter100|18300_ , \new_Sorter100|18399_ , \new_Sorter100|18301_ ,
    \new_Sorter100|18302_ , \new_Sorter100|18303_ , \new_Sorter100|18304_ ,
    \new_Sorter100|18305_ , \new_Sorter100|18306_ , \new_Sorter100|18307_ ,
    \new_Sorter100|18308_ , \new_Sorter100|18309_ , \new_Sorter100|18310_ ,
    \new_Sorter100|18311_ , \new_Sorter100|18312_ , \new_Sorter100|18313_ ,
    \new_Sorter100|18314_ , \new_Sorter100|18315_ , \new_Sorter100|18316_ ,
    \new_Sorter100|18317_ , \new_Sorter100|18318_ , \new_Sorter100|18319_ ,
    \new_Sorter100|18320_ , \new_Sorter100|18321_ , \new_Sorter100|18322_ ,
    \new_Sorter100|18323_ , \new_Sorter100|18324_ , \new_Sorter100|18325_ ,
    \new_Sorter100|18326_ , \new_Sorter100|18327_ , \new_Sorter100|18328_ ,
    \new_Sorter100|18329_ , \new_Sorter100|18330_ , \new_Sorter100|18331_ ,
    \new_Sorter100|18332_ , \new_Sorter100|18333_ , \new_Sorter100|18334_ ,
    \new_Sorter100|18335_ , \new_Sorter100|18336_ , \new_Sorter100|18337_ ,
    \new_Sorter100|18338_ , \new_Sorter100|18339_ , \new_Sorter100|18340_ ,
    \new_Sorter100|18341_ , \new_Sorter100|18342_ , \new_Sorter100|18343_ ,
    \new_Sorter100|18344_ , \new_Sorter100|18345_ , \new_Sorter100|18346_ ,
    \new_Sorter100|18347_ , \new_Sorter100|18348_ , \new_Sorter100|18349_ ,
    \new_Sorter100|18350_ , \new_Sorter100|18351_ , \new_Sorter100|18352_ ,
    \new_Sorter100|18353_ , \new_Sorter100|18354_ , \new_Sorter100|18355_ ,
    \new_Sorter100|18356_ , \new_Sorter100|18357_ , \new_Sorter100|18358_ ,
    \new_Sorter100|18359_ , \new_Sorter100|18360_ , \new_Sorter100|18361_ ,
    \new_Sorter100|18362_ , \new_Sorter100|18363_ , \new_Sorter100|18364_ ,
    \new_Sorter100|18365_ , \new_Sorter100|18366_ , \new_Sorter100|18367_ ,
    \new_Sorter100|18368_ , \new_Sorter100|18369_ , \new_Sorter100|18370_ ,
    \new_Sorter100|18371_ , \new_Sorter100|18372_ , \new_Sorter100|18373_ ,
    \new_Sorter100|18374_ , \new_Sorter100|18375_ , \new_Sorter100|18376_ ,
    \new_Sorter100|18377_ , \new_Sorter100|18378_ , \new_Sorter100|18379_ ,
    \new_Sorter100|18380_ , \new_Sorter100|18381_ , \new_Sorter100|18382_ ,
    \new_Sorter100|18383_ , \new_Sorter100|18384_ , \new_Sorter100|18385_ ,
    \new_Sorter100|18386_ , \new_Sorter100|18387_ , \new_Sorter100|18388_ ,
    \new_Sorter100|18389_ , \new_Sorter100|18390_ , \new_Sorter100|18391_ ,
    \new_Sorter100|18392_ , \new_Sorter100|18393_ , \new_Sorter100|18394_ ,
    \new_Sorter100|18395_ , \new_Sorter100|18396_ , \new_Sorter100|18397_ ,
    \new_Sorter100|18398_ , \new_Sorter100|18400_ , \new_Sorter100|18401_ ,
    \new_Sorter100|18402_ , \new_Sorter100|18403_ , \new_Sorter100|18404_ ,
    \new_Sorter100|18405_ , \new_Sorter100|18406_ , \new_Sorter100|18407_ ,
    \new_Sorter100|18408_ , \new_Sorter100|18409_ , \new_Sorter100|18410_ ,
    \new_Sorter100|18411_ , \new_Sorter100|18412_ , \new_Sorter100|18413_ ,
    \new_Sorter100|18414_ , \new_Sorter100|18415_ , \new_Sorter100|18416_ ,
    \new_Sorter100|18417_ , \new_Sorter100|18418_ , \new_Sorter100|18419_ ,
    \new_Sorter100|18420_ , \new_Sorter100|18421_ , \new_Sorter100|18422_ ,
    \new_Sorter100|18423_ , \new_Sorter100|18424_ , \new_Sorter100|18425_ ,
    \new_Sorter100|18426_ , \new_Sorter100|18427_ , \new_Sorter100|18428_ ,
    \new_Sorter100|18429_ , \new_Sorter100|18430_ , \new_Sorter100|18431_ ,
    \new_Sorter100|18432_ , \new_Sorter100|18433_ , \new_Sorter100|18434_ ,
    \new_Sorter100|18435_ , \new_Sorter100|18436_ , \new_Sorter100|18437_ ,
    \new_Sorter100|18438_ , \new_Sorter100|18439_ , \new_Sorter100|18440_ ,
    \new_Sorter100|18441_ , \new_Sorter100|18442_ , \new_Sorter100|18443_ ,
    \new_Sorter100|18444_ , \new_Sorter100|18445_ , \new_Sorter100|18446_ ,
    \new_Sorter100|18447_ , \new_Sorter100|18448_ , \new_Sorter100|18449_ ,
    \new_Sorter100|18450_ , \new_Sorter100|18451_ , \new_Sorter100|18452_ ,
    \new_Sorter100|18453_ , \new_Sorter100|18454_ , \new_Sorter100|18455_ ,
    \new_Sorter100|18456_ , \new_Sorter100|18457_ , \new_Sorter100|18458_ ,
    \new_Sorter100|18459_ , \new_Sorter100|18460_ , \new_Sorter100|18461_ ,
    \new_Sorter100|18462_ , \new_Sorter100|18463_ , \new_Sorter100|18464_ ,
    \new_Sorter100|18465_ , \new_Sorter100|18466_ , \new_Sorter100|18467_ ,
    \new_Sorter100|18468_ , \new_Sorter100|18469_ , \new_Sorter100|18470_ ,
    \new_Sorter100|18471_ , \new_Sorter100|18472_ , \new_Sorter100|18473_ ,
    \new_Sorter100|18474_ , \new_Sorter100|18475_ , \new_Sorter100|18476_ ,
    \new_Sorter100|18477_ , \new_Sorter100|18478_ , \new_Sorter100|18479_ ,
    \new_Sorter100|18480_ , \new_Sorter100|18481_ , \new_Sorter100|18482_ ,
    \new_Sorter100|18483_ , \new_Sorter100|18484_ , \new_Sorter100|18485_ ,
    \new_Sorter100|18486_ , \new_Sorter100|18487_ , \new_Sorter100|18488_ ,
    \new_Sorter100|18489_ , \new_Sorter100|18490_ , \new_Sorter100|18491_ ,
    \new_Sorter100|18492_ , \new_Sorter100|18493_ , \new_Sorter100|18494_ ,
    \new_Sorter100|18495_ , \new_Sorter100|18496_ , \new_Sorter100|18497_ ,
    \new_Sorter100|18498_ , \new_Sorter100|18499_ , \new_Sorter100|18500_ ,
    \new_Sorter100|18599_ , \new_Sorter100|18501_ , \new_Sorter100|18502_ ,
    \new_Sorter100|18503_ , \new_Sorter100|18504_ , \new_Sorter100|18505_ ,
    \new_Sorter100|18506_ , \new_Sorter100|18507_ , \new_Sorter100|18508_ ,
    \new_Sorter100|18509_ , \new_Sorter100|18510_ , \new_Sorter100|18511_ ,
    \new_Sorter100|18512_ , \new_Sorter100|18513_ , \new_Sorter100|18514_ ,
    \new_Sorter100|18515_ , \new_Sorter100|18516_ , \new_Sorter100|18517_ ,
    \new_Sorter100|18518_ , \new_Sorter100|18519_ , \new_Sorter100|18520_ ,
    \new_Sorter100|18521_ , \new_Sorter100|18522_ , \new_Sorter100|18523_ ,
    \new_Sorter100|18524_ , \new_Sorter100|18525_ , \new_Sorter100|18526_ ,
    \new_Sorter100|18527_ , \new_Sorter100|18528_ , \new_Sorter100|18529_ ,
    \new_Sorter100|18530_ , \new_Sorter100|18531_ , \new_Sorter100|18532_ ,
    \new_Sorter100|18533_ , \new_Sorter100|18534_ , \new_Sorter100|18535_ ,
    \new_Sorter100|18536_ , \new_Sorter100|18537_ , \new_Sorter100|18538_ ,
    \new_Sorter100|18539_ , \new_Sorter100|18540_ , \new_Sorter100|18541_ ,
    \new_Sorter100|18542_ , \new_Sorter100|18543_ , \new_Sorter100|18544_ ,
    \new_Sorter100|18545_ , \new_Sorter100|18546_ , \new_Sorter100|18547_ ,
    \new_Sorter100|18548_ , \new_Sorter100|18549_ , \new_Sorter100|18550_ ,
    \new_Sorter100|18551_ , \new_Sorter100|18552_ , \new_Sorter100|18553_ ,
    \new_Sorter100|18554_ , \new_Sorter100|18555_ , \new_Sorter100|18556_ ,
    \new_Sorter100|18557_ , \new_Sorter100|18558_ , \new_Sorter100|18559_ ,
    \new_Sorter100|18560_ , \new_Sorter100|18561_ , \new_Sorter100|18562_ ,
    \new_Sorter100|18563_ , \new_Sorter100|18564_ , \new_Sorter100|18565_ ,
    \new_Sorter100|18566_ , \new_Sorter100|18567_ , \new_Sorter100|18568_ ,
    \new_Sorter100|18569_ , \new_Sorter100|18570_ , \new_Sorter100|18571_ ,
    \new_Sorter100|18572_ , \new_Sorter100|18573_ , \new_Sorter100|18574_ ,
    \new_Sorter100|18575_ , \new_Sorter100|18576_ , \new_Sorter100|18577_ ,
    \new_Sorter100|18578_ , \new_Sorter100|18579_ , \new_Sorter100|18580_ ,
    \new_Sorter100|18581_ , \new_Sorter100|18582_ , \new_Sorter100|18583_ ,
    \new_Sorter100|18584_ , \new_Sorter100|18585_ , \new_Sorter100|18586_ ,
    \new_Sorter100|18587_ , \new_Sorter100|18588_ , \new_Sorter100|18589_ ,
    \new_Sorter100|18590_ , \new_Sorter100|18591_ , \new_Sorter100|18592_ ,
    \new_Sorter100|18593_ , \new_Sorter100|18594_ , \new_Sorter100|18595_ ,
    \new_Sorter100|18596_ , \new_Sorter100|18597_ , \new_Sorter100|18598_ ,
    \new_Sorter100|18600_ , \new_Sorter100|18601_ , \new_Sorter100|18602_ ,
    \new_Sorter100|18603_ , \new_Sorter100|18604_ , \new_Sorter100|18605_ ,
    \new_Sorter100|18606_ , \new_Sorter100|18607_ , \new_Sorter100|18608_ ,
    \new_Sorter100|18609_ , \new_Sorter100|18610_ , \new_Sorter100|18611_ ,
    \new_Sorter100|18612_ , \new_Sorter100|18613_ , \new_Sorter100|18614_ ,
    \new_Sorter100|18615_ , \new_Sorter100|18616_ , \new_Sorter100|18617_ ,
    \new_Sorter100|18618_ , \new_Sorter100|18619_ , \new_Sorter100|18620_ ,
    \new_Sorter100|18621_ , \new_Sorter100|18622_ , \new_Sorter100|18623_ ,
    \new_Sorter100|18624_ , \new_Sorter100|18625_ , \new_Sorter100|18626_ ,
    \new_Sorter100|18627_ , \new_Sorter100|18628_ , \new_Sorter100|18629_ ,
    \new_Sorter100|18630_ , \new_Sorter100|18631_ , \new_Sorter100|18632_ ,
    \new_Sorter100|18633_ , \new_Sorter100|18634_ , \new_Sorter100|18635_ ,
    \new_Sorter100|18636_ , \new_Sorter100|18637_ , \new_Sorter100|18638_ ,
    \new_Sorter100|18639_ , \new_Sorter100|18640_ , \new_Sorter100|18641_ ,
    \new_Sorter100|18642_ , \new_Sorter100|18643_ , \new_Sorter100|18644_ ,
    \new_Sorter100|18645_ , \new_Sorter100|18646_ , \new_Sorter100|18647_ ,
    \new_Sorter100|18648_ , \new_Sorter100|18649_ , \new_Sorter100|18650_ ,
    \new_Sorter100|18651_ , \new_Sorter100|18652_ , \new_Sorter100|18653_ ,
    \new_Sorter100|18654_ , \new_Sorter100|18655_ , \new_Sorter100|18656_ ,
    \new_Sorter100|18657_ , \new_Sorter100|18658_ , \new_Sorter100|18659_ ,
    \new_Sorter100|18660_ , \new_Sorter100|18661_ , \new_Sorter100|18662_ ,
    \new_Sorter100|18663_ , \new_Sorter100|18664_ , \new_Sorter100|18665_ ,
    \new_Sorter100|18666_ , \new_Sorter100|18667_ , \new_Sorter100|18668_ ,
    \new_Sorter100|18669_ , \new_Sorter100|18670_ , \new_Sorter100|18671_ ,
    \new_Sorter100|18672_ , \new_Sorter100|18673_ , \new_Sorter100|18674_ ,
    \new_Sorter100|18675_ , \new_Sorter100|18676_ , \new_Sorter100|18677_ ,
    \new_Sorter100|18678_ , \new_Sorter100|18679_ , \new_Sorter100|18680_ ,
    \new_Sorter100|18681_ , \new_Sorter100|18682_ , \new_Sorter100|18683_ ,
    \new_Sorter100|18684_ , \new_Sorter100|18685_ , \new_Sorter100|18686_ ,
    \new_Sorter100|18687_ , \new_Sorter100|18688_ , \new_Sorter100|18689_ ,
    \new_Sorter100|18690_ , \new_Sorter100|18691_ , \new_Sorter100|18692_ ,
    \new_Sorter100|18693_ , \new_Sorter100|18694_ , \new_Sorter100|18695_ ,
    \new_Sorter100|18696_ , \new_Sorter100|18697_ , \new_Sorter100|18698_ ,
    \new_Sorter100|18699_ , \new_Sorter100|18700_ , \new_Sorter100|18799_ ,
    \new_Sorter100|18701_ , \new_Sorter100|18702_ , \new_Sorter100|18703_ ,
    \new_Sorter100|18704_ , \new_Sorter100|18705_ , \new_Sorter100|18706_ ,
    \new_Sorter100|18707_ , \new_Sorter100|18708_ , \new_Sorter100|18709_ ,
    \new_Sorter100|18710_ , \new_Sorter100|18711_ , \new_Sorter100|18712_ ,
    \new_Sorter100|18713_ , \new_Sorter100|18714_ , \new_Sorter100|18715_ ,
    \new_Sorter100|18716_ , \new_Sorter100|18717_ , \new_Sorter100|18718_ ,
    \new_Sorter100|18719_ , \new_Sorter100|18720_ , \new_Sorter100|18721_ ,
    \new_Sorter100|18722_ , \new_Sorter100|18723_ , \new_Sorter100|18724_ ,
    \new_Sorter100|18725_ , \new_Sorter100|18726_ , \new_Sorter100|18727_ ,
    \new_Sorter100|18728_ , \new_Sorter100|18729_ , \new_Sorter100|18730_ ,
    \new_Sorter100|18731_ , \new_Sorter100|18732_ , \new_Sorter100|18733_ ,
    \new_Sorter100|18734_ , \new_Sorter100|18735_ , \new_Sorter100|18736_ ,
    \new_Sorter100|18737_ , \new_Sorter100|18738_ , \new_Sorter100|18739_ ,
    \new_Sorter100|18740_ , \new_Sorter100|18741_ , \new_Sorter100|18742_ ,
    \new_Sorter100|18743_ , \new_Sorter100|18744_ , \new_Sorter100|18745_ ,
    \new_Sorter100|18746_ , \new_Sorter100|18747_ , \new_Sorter100|18748_ ,
    \new_Sorter100|18749_ , \new_Sorter100|18750_ , \new_Sorter100|18751_ ,
    \new_Sorter100|18752_ , \new_Sorter100|18753_ , \new_Sorter100|18754_ ,
    \new_Sorter100|18755_ , \new_Sorter100|18756_ , \new_Sorter100|18757_ ,
    \new_Sorter100|18758_ , \new_Sorter100|18759_ , \new_Sorter100|18760_ ,
    \new_Sorter100|18761_ , \new_Sorter100|18762_ , \new_Sorter100|18763_ ,
    \new_Sorter100|18764_ , \new_Sorter100|18765_ , \new_Sorter100|18766_ ,
    \new_Sorter100|18767_ , \new_Sorter100|18768_ , \new_Sorter100|18769_ ,
    \new_Sorter100|18770_ , \new_Sorter100|18771_ , \new_Sorter100|18772_ ,
    \new_Sorter100|18773_ , \new_Sorter100|18774_ , \new_Sorter100|18775_ ,
    \new_Sorter100|18776_ , \new_Sorter100|18777_ , \new_Sorter100|18778_ ,
    \new_Sorter100|18779_ , \new_Sorter100|18780_ , \new_Sorter100|18781_ ,
    \new_Sorter100|18782_ , \new_Sorter100|18783_ , \new_Sorter100|18784_ ,
    \new_Sorter100|18785_ , \new_Sorter100|18786_ , \new_Sorter100|18787_ ,
    \new_Sorter100|18788_ , \new_Sorter100|18789_ , \new_Sorter100|18790_ ,
    \new_Sorter100|18791_ , \new_Sorter100|18792_ , \new_Sorter100|18793_ ,
    \new_Sorter100|18794_ , \new_Sorter100|18795_ , \new_Sorter100|18796_ ,
    \new_Sorter100|18797_ , \new_Sorter100|18798_ , \new_Sorter100|18800_ ,
    \new_Sorter100|18801_ , \new_Sorter100|18802_ , \new_Sorter100|18803_ ,
    \new_Sorter100|18804_ , \new_Sorter100|18805_ , \new_Sorter100|18806_ ,
    \new_Sorter100|18807_ , \new_Sorter100|18808_ , \new_Sorter100|18809_ ,
    \new_Sorter100|18810_ , \new_Sorter100|18811_ , \new_Sorter100|18812_ ,
    \new_Sorter100|18813_ , \new_Sorter100|18814_ , \new_Sorter100|18815_ ,
    \new_Sorter100|18816_ , \new_Sorter100|18817_ , \new_Sorter100|18818_ ,
    \new_Sorter100|18819_ , \new_Sorter100|18820_ , \new_Sorter100|18821_ ,
    \new_Sorter100|18822_ , \new_Sorter100|18823_ , \new_Sorter100|18824_ ,
    \new_Sorter100|18825_ , \new_Sorter100|18826_ , \new_Sorter100|18827_ ,
    \new_Sorter100|18828_ , \new_Sorter100|18829_ , \new_Sorter100|18830_ ,
    \new_Sorter100|18831_ , \new_Sorter100|18832_ , \new_Sorter100|18833_ ,
    \new_Sorter100|18834_ , \new_Sorter100|18835_ , \new_Sorter100|18836_ ,
    \new_Sorter100|18837_ , \new_Sorter100|18838_ , \new_Sorter100|18839_ ,
    \new_Sorter100|18840_ , \new_Sorter100|18841_ , \new_Sorter100|18842_ ,
    \new_Sorter100|18843_ , \new_Sorter100|18844_ , \new_Sorter100|18845_ ,
    \new_Sorter100|18846_ , \new_Sorter100|18847_ , \new_Sorter100|18848_ ,
    \new_Sorter100|18849_ , \new_Sorter100|18850_ , \new_Sorter100|18851_ ,
    \new_Sorter100|18852_ , \new_Sorter100|18853_ , \new_Sorter100|18854_ ,
    \new_Sorter100|18855_ , \new_Sorter100|18856_ , \new_Sorter100|18857_ ,
    \new_Sorter100|18858_ , \new_Sorter100|18859_ , \new_Sorter100|18860_ ,
    \new_Sorter100|18861_ , \new_Sorter100|18862_ , \new_Sorter100|18863_ ,
    \new_Sorter100|18864_ , \new_Sorter100|18865_ , \new_Sorter100|18866_ ,
    \new_Sorter100|18867_ , \new_Sorter100|18868_ , \new_Sorter100|18869_ ,
    \new_Sorter100|18870_ , \new_Sorter100|18871_ , \new_Sorter100|18872_ ,
    \new_Sorter100|18873_ , \new_Sorter100|18874_ , \new_Sorter100|18875_ ,
    \new_Sorter100|18876_ , \new_Sorter100|18877_ , \new_Sorter100|18878_ ,
    \new_Sorter100|18879_ , \new_Sorter100|18880_ , \new_Sorter100|18881_ ,
    \new_Sorter100|18882_ , \new_Sorter100|18883_ , \new_Sorter100|18884_ ,
    \new_Sorter100|18885_ , \new_Sorter100|18886_ , \new_Sorter100|18887_ ,
    \new_Sorter100|18888_ , \new_Sorter100|18889_ , \new_Sorter100|18890_ ,
    \new_Sorter100|18891_ , \new_Sorter100|18892_ , \new_Sorter100|18893_ ,
    \new_Sorter100|18894_ , \new_Sorter100|18895_ , \new_Sorter100|18896_ ,
    \new_Sorter100|18897_ , \new_Sorter100|18898_ , \new_Sorter100|18899_ ,
    \new_Sorter100|18900_ , \new_Sorter100|18999_ , \new_Sorter100|18901_ ,
    \new_Sorter100|18902_ , \new_Sorter100|18903_ , \new_Sorter100|18904_ ,
    \new_Sorter100|18905_ , \new_Sorter100|18906_ , \new_Sorter100|18907_ ,
    \new_Sorter100|18908_ , \new_Sorter100|18909_ , \new_Sorter100|18910_ ,
    \new_Sorter100|18911_ , \new_Sorter100|18912_ , \new_Sorter100|18913_ ,
    \new_Sorter100|18914_ , \new_Sorter100|18915_ , \new_Sorter100|18916_ ,
    \new_Sorter100|18917_ , \new_Sorter100|18918_ , \new_Sorter100|18919_ ,
    \new_Sorter100|18920_ , \new_Sorter100|18921_ , \new_Sorter100|18922_ ,
    \new_Sorter100|18923_ , \new_Sorter100|18924_ , \new_Sorter100|18925_ ,
    \new_Sorter100|18926_ , \new_Sorter100|18927_ , \new_Sorter100|18928_ ,
    \new_Sorter100|18929_ , \new_Sorter100|18930_ , \new_Sorter100|18931_ ,
    \new_Sorter100|18932_ , \new_Sorter100|18933_ , \new_Sorter100|18934_ ,
    \new_Sorter100|18935_ , \new_Sorter100|18936_ , \new_Sorter100|18937_ ,
    \new_Sorter100|18938_ , \new_Sorter100|18939_ , \new_Sorter100|18940_ ,
    \new_Sorter100|18941_ , \new_Sorter100|18942_ , \new_Sorter100|18943_ ,
    \new_Sorter100|18944_ , \new_Sorter100|18945_ , \new_Sorter100|18946_ ,
    \new_Sorter100|18947_ , \new_Sorter100|18948_ , \new_Sorter100|18949_ ,
    \new_Sorter100|18950_ , \new_Sorter100|18951_ , \new_Sorter100|18952_ ,
    \new_Sorter100|18953_ , \new_Sorter100|18954_ , \new_Sorter100|18955_ ,
    \new_Sorter100|18956_ , \new_Sorter100|18957_ , \new_Sorter100|18958_ ,
    \new_Sorter100|18959_ , \new_Sorter100|18960_ , \new_Sorter100|18961_ ,
    \new_Sorter100|18962_ , \new_Sorter100|18963_ , \new_Sorter100|18964_ ,
    \new_Sorter100|18965_ , \new_Sorter100|18966_ , \new_Sorter100|18967_ ,
    \new_Sorter100|18968_ , \new_Sorter100|18969_ , \new_Sorter100|18970_ ,
    \new_Sorter100|18971_ , \new_Sorter100|18972_ , \new_Sorter100|18973_ ,
    \new_Sorter100|18974_ , \new_Sorter100|18975_ , \new_Sorter100|18976_ ,
    \new_Sorter100|18977_ , \new_Sorter100|18978_ , \new_Sorter100|18979_ ,
    \new_Sorter100|18980_ , \new_Sorter100|18981_ , \new_Sorter100|18982_ ,
    \new_Sorter100|18983_ , \new_Sorter100|18984_ , \new_Sorter100|18985_ ,
    \new_Sorter100|18986_ , \new_Sorter100|18987_ , \new_Sorter100|18988_ ,
    \new_Sorter100|18989_ , \new_Sorter100|18990_ , \new_Sorter100|18991_ ,
    \new_Sorter100|18992_ , \new_Sorter100|18993_ , \new_Sorter100|18994_ ,
    \new_Sorter100|18995_ , \new_Sorter100|18996_ , \new_Sorter100|18997_ ,
    \new_Sorter100|18998_ , \new_Sorter100|19000_ , \new_Sorter100|19001_ ,
    \new_Sorter100|19002_ , \new_Sorter100|19003_ , \new_Sorter100|19004_ ,
    \new_Sorter100|19005_ , \new_Sorter100|19006_ , \new_Sorter100|19007_ ,
    \new_Sorter100|19008_ , \new_Sorter100|19009_ , \new_Sorter100|19010_ ,
    \new_Sorter100|19011_ , \new_Sorter100|19012_ , \new_Sorter100|19013_ ,
    \new_Sorter100|19014_ , \new_Sorter100|19015_ , \new_Sorter100|19016_ ,
    \new_Sorter100|19017_ , \new_Sorter100|19018_ , \new_Sorter100|19019_ ,
    \new_Sorter100|19020_ , \new_Sorter100|19021_ , \new_Sorter100|19022_ ,
    \new_Sorter100|19023_ , \new_Sorter100|19024_ , \new_Sorter100|19025_ ,
    \new_Sorter100|19026_ , \new_Sorter100|19027_ , \new_Sorter100|19028_ ,
    \new_Sorter100|19029_ , \new_Sorter100|19030_ , \new_Sorter100|19031_ ,
    \new_Sorter100|19032_ , \new_Sorter100|19033_ , \new_Sorter100|19034_ ,
    \new_Sorter100|19035_ , \new_Sorter100|19036_ , \new_Sorter100|19037_ ,
    \new_Sorter100|19038_ , \new_Sorter100|19039_ , \new_Sorter100|19040_ ,
    \new_Sorter100|19041_ , \new_Sorter100|19042_ , \new_Sorter100|19043_ ,
    \new_Sorter100|19044_ , \new_Sorter100|19045_ , \new_Sorter100|19046_ ,
    \new_Sorter100|19047_ , \new_Sorter100|19048_ , \new_Sorter100|19049_ ,
    \new_Sorter100|19050_ , \new_Sorter100|19051_ , \new_Sorter100|19052_ ,
    \new_Sorter100|19053_ , \new_Sorter100|19054_ , \new_Sorter100|19055_ ,
    \new_Sorter100|19056_ , \new_Sorter100|19057_ , \new_Sorter100|19058_ ,
    \new_Sorter100|19059_ , \new_Sorter100|19060_ , \new_Sorter100|19061_ ,
    \new_Sorter100|19062_ , \new_Sorter100|19063_ , \new_Sorter100|19064_ ,
    \new_Sorter100|19065_ , \new_Sorter100|19066_ , \new_Sorter100|19067_ ,
    \new_Sorter100|19068_ , \new_Sorter100|19069_ , \new_Sorter100|19070_ ,
    \new_Sorter100|19071_ , \new_Sorter100|19072_ , \new_Sorter100|19073_ ,
    \new_Sorter100|19074_ , \new_Sorter100|19075_ , \new_Sorter100|19076_ ,
    \new_Sorter100|19077_ , \new_Sorter100|19078_ , \new_Sorter100|19079_ ,
    \new_Sorter100|19080_ , \new_Sorter100|19081_ , \new_Sorter100|19082_ ,
    \new_Sorter100|19083_ , \new_Sorter100|19084_ , \new_Sorter100|19085_ ,
    \new_Sorter100|19086_ , \new_Sorter100|19087_ , \new_Sorter100|19088_ ,
    \new_Sorter100|19089_ , \new_Sorter100|19090_ , \new_Sorter100|19091_ ,
    \new_Sorter100|19092_ , \new_Sorter100|19093_ , \new_Sorter100|19094_ ,
    \new_Sorter100|19095_ , \new_Sorter100|19096_ , \new_Sorter100|19097_ ,
    \new_Sorter100|19098_ , \new_Sorter100|19099_ , \new_Sorter100|19100_ ,
    \new_Sorter100|19199_ , \new_Sorter100|19101_ , \new_Sorter100|19102_ ,
    \new_Sorter100|19103_ , \new_Sorter100|19104_ , \new_Sorter100|19105_ ,
    \new_Sorter100|19106_ , \new_Sorter100|19107_ , \new_Sorter100|19108_ ,
    \new_Sorter100|19109_ , \new_Sorter100|19110_ , \new_Sorter100|19111_ ,
    \new_Sorter100|19112_ , \new_Sorter100|19113_ , \new_Sorter100|19114_ ,
    \new_Sorter100|19115_ , \new_Sorter100|19116_ , \new_Sorter100|19117_ ,
    \new_Sorter100|19118_ , \new_Sorter100|19119_ , \new_Sorter100|19120_ ,
    \new_Sorter100|19121_ , \new_Sorter100|19122_ , \new_Sorter100|19123_ ,
    \new_Sorter100|19124_ , \new_Sorter100|19125_ , \new_Sorter100|19126_ ,
    \new_Sorter100|19127_ , \new_Sorter100|19128_ , \new_Sorter100|19129_ ,
    \new_Sorter100|19130_ , \new_Sorter100|19131_ , \new_Sorter100|19132_ ,
    \new_Sorter100|19133_ , \new_Sorter100|19134_ , \new_Sorter100|19135_ ,
    \new_Sorter100|19136_ , \new_Sorter100|19137_ , \new_Sorter100|19138_ ,
    \new_Sorter100|19139_ , \new_Sorter100|19140_ , \new_Sorter100|19141_ ,
    \new_Sorter100|19142_ , \new_Sorter100|19143_ , \new_Sorter100|19144_ ,
    \new_Sorter100|19145_ , \new_Sorter100|19146_ , \new_Sorter100|19147_ ,
    \new_Sorter100|19148_ , \new_Sorter100|19149_ , \new_Sorter100|19150_ ,
    \new_Sorter100|19151_ , \new_Sorter100|19152_ , \new_Sorter100|19153_ ,
    \new_Sorter100|19154_ , \new_Sorter100|19155_ , \new_Sorter100|19156_ ,
    \new_Sorter100|19157_ , \new_Sorter100|19158_ , \new_Sorter100|19159_ ,
    \new_Sorter100|19160_ , \new_Sorter100|19161_ , \new_Sorter100|19162_ ,
    \new_Sorter100|19163_ , \new_Sorter100|19164_ , \new_Sorter100|19165_ ,
    \new_Sorter100|19166_ , \new_Sorter100|19167_ , \new_Sorter100|19168_ ,
    \new_Sorter100|19169_ , \new_Sorter100|19170_ , \new_Sorter100|19171_ ,
    \new_Sorter100|19172_ , \new_Sorter100|19173_ , \new_Sorter100|19174_ ,
    \new_Sorter100|19175_ , \new_Sorter100|19176_ , \new_Sorter100|19177_ ,
    \new_Sorter100|19178_ , \new_Sorter100|19179_ , \new_Sorter100|19180_ ,
    \new_Sorter100|19181_ , \new_Sorter100|19182_ , \new_Sorter100|19183_ ,
    \new_Sorter100|19184_ , \new_Sorter100|19185_ , \new_Sorter100|19186_ ,
    \new_Sorter100|19187_ , \new_Sorter100|19188_ , \new_Sorter100|19189_ ,
    \new_Sorter100|19190_ , \new_Sorter100|19191_ , \new_Sorter100|19192_ ,
    \new_Sorter100|19193_ , \new_Sorter100|19194_ , \new_Sorter100|19195_ ,
    \new_Sorter100|19196_ , \new_Sorter100|19197_ , \new_Sorter100|19198_ ,
    \new_Sorter100|19200_ , \new_Sorter100|19201_ , \new_Sorter100|19202_ ,
    \new_Sorter100|19203_ , \new_Sorter100|19204_ , \new_Sorter100|19205_ ,
    \new_Sorter100|19206_ , \new_Sorter100|19207_ , \new_Sorter100|19208_ ,
    \new_Sorter100|19209_ , \new_Sorter100|19210_ , \new_Sorter100|19211_ ,
    \new_Sorter100|19212_ , \new_Sorter100|19213_ , \new_Sorter100|19214_ ,
    \new_Sorter100|19215_ , \new_Sorter100|19216_ , \new_Sorter100|19217_ ,
    \new_Sorter100|19218_ , \new_Sorter100|19219_ , \new_Sorter100|19220_ ,
    \new_Sorter100|19221_ , \new_Sorter100|19222_ , \new_Sorter100|19223_ ,
    \new_Sorter100|19224_ , \new_Sorter100|19225_ , \new_Sorter100|19226_ ,
    \new_Sorter100|19227_ , \new_Sorter100|19228_ , \new_Sorter100|19229_ ,
    \new_Sorter100|19230_ , \new_Sorter100|19231_ , \new_Sorter100|19232_ ,
    \new_Sorter100|19233_ , \new_Sorter100|19234_ , \new_Sorter100|19235_ ,
    \new_Sorter100|19236_ , \new_Sorter100|19237_ , \new_Sorter100|19238_ ,
    \new_Sorter100|19239_ , \new_Sorter100|19240_ , \new_Sorter100|19241_ ,
    \new_Sorter100|19242_ , \new_Sorter100|19243_ , \new_Sorter100|19244_ ,
    \new_Sorter100|19245_ , \new_Sorter100|19246_ , \new_Sorter100|19247_ ,
    \new_Sorter100|19248_ , \new_Sorter100|19249_ , \new_Sorter100|19250_ ,
    \new_Sorter100|19251_ , \new_Sorter100|19252_ , \new_Sorter100|19253_ ,
    \new_Sorter100|19254_ , \new_Sorter100|19255_ , \new_Sorter100|19256_ ,
    \new_Sorter100|19257_ , \new_Sorter100|19258_ , \new_Sorter100|19259_ ,
    \new_Sorter100|19260_ , \new_Sorter100|19261_ , \new_Sorter100|19262_ ,
    \new_Sorter100|19263_ , \new_Sorter100|19264_ , \new_Sorter100|19265_ ,
    \new_Sorter100|19266_ , \new_Sorter100|19267_ , \new_Sorter100|19268_ ,
    \new_Sorter100|19269_ , \new_Sorter100|19270_ , \new_Sorter100|19271_ ,
    \new_Sorter100|19272_ , \new_Sorter100|19273_ , \new_Sorter100|19274_ ,
    \new_Sorter100|19275_ , \new_Sorter100|19276_ , \new_Sorter100|19277_ ,
    \new_Sorter100|19278_ , \new_Sorter100|19279_ , \new_Sorter100|19280_ ,
    \new_Sorter100|19281_ , \new_Sorter100|19282_ , \new_Sorter100|19283_ ,
    \new_Sorter100|19284_ , \new_Sorter100|19285_ , \new_Sorter100|19286_ ,
    \new_Sorter100|19287_ , \new_Sorter100|19288_ , \new_Sorter100|19289_ ,
    \new_Sorter100|19290_ , \new_Sorter100|19291_ , \new_Sorter100|19292_ ,
    \new_Sorter100|19293_ , \new_Sorter100|19294_ , \new_Sorter100|19295_ ,
    \new_Sorter100|19296_ , \new_Sorter100|19297_ , \new_Sorter100|19298_ ,
    \new_Sorter100|19299_ , \new_Sorter100|19300_ , \new_Sorter100|19399_ ,
    \new_Sorter100|19301_ , \new_Sorter100|19302_ , \new_Sorter100|19303_ ,
    \new_Sorter100|19304_ , \new_Sorter100|19305_ , \new_Sorter100|19306_ ,
    \new_Sorter100|19307_ , \new_Sorter100|19308_ , \new_Sorter100|19309_ ,
    \new_Sorter100|19310_ , \new_Sorter100|19311_ , \new_Sorter100|19312_ ,
    \new_Sorter100|19313_ , \new_Sorter100|19314_ , \new_Sorter100|19315_ ,
    \new_Sorter100|19316_ , \new_Sorter100|19317_ , \new_Sorter100|19318_ ,
    \new_Sorter100|19319_ , \new_Sorter100|19320_ , \new_Sorter100|19321_ ,
    \new_Sorter100|19322_ , \new_Sorter100|19323_ , \new_Sorter100|19324_ ,
    \new_Sorter100|19325_ , \new_Sorter100|19326_ , \new_Sorter100|19327_ ,
    \new_Sorter100|19328_ , \new_Sorter100|19329_ , \new_Sorter100|19330_ ,
    \new_Sorter100|19331_ , \new_Sorter100|19332_ , \new_Sorter100|19333_ ,
    \new_Sorter100|19334_ , \new_Sorter100|19335_ , \new_Sorter100|19336_ ,
    \new_Sorter100|19337_ , \new_Sorter100|19338_ , \new_Sorter100|19339_ ,
    \new_Sorter100|19340_ , \new_Sorter100|19341_ , \new_Sorter100|19342_ ,
    \new_Sorter100|19343_ , \new_Sorter100|19344_ , \new_Sorter100|19345_ ,
    \new_Sorter100|19346_ , \new_Sorter100|19347_ , \new_Sorter100|19348_ ,
    \new_Sorter100|19349_ , \new_Sorter100|19350_ , \new_Sorter100|19351_ ,
    \new_Sorter100|19352_ , \new_Sorter100|19353_ , \new_Sorter100|19354_ ,
    \new_Sorter100|19355_ , \new_Sorter100|19356_ , \new_Sorter100|19357_ ,
    \new_Sorter100|19358_ , \new_Sorter100|19359_ , \new_Sorter100|19360_ ,
    \new_Sorter100|19361_ , \new_Sorter100|19362_ , \new_Sorter100|19363_ ,
    \new_Sorter100|19364_ , \new_Sorter100|19365_ , \new_Sorter100|19366_ ,
    \new_Sorter100|19367_ , \new_Sorter100|19368_ , \new_Sorter100|19369_ ,
    \new_Sorter100|19370_ , \new_Sorter100|19371_ , \new_Sorter100|19372_ ,
    \new_Sorter100|19373_ , \new_Sorter100|19374_ , \new_Sorter100|19375_ ,
    \new_Sorter100|19376_ , \new_Sorter100|19377_ , \new_Sorter100|19378_ ,
    \new_Sorter100|19379_ , \new_Sorter100|19380_ , \new_Sorter100|19381_ ,
    \new_Sorter100|19382_ , \new_Sorter100|19383_ , \new_Sorter100|19384_ ,
    \new_Sorter100|19385_ , \new_Sorter100|19386_ , \new_Sorter100|19387_ ,
    \new_Sorter100|19388_ , \new_Sorter100|19389_ , \new_Sorter100|19390_ ,
    \new_Sorter100|19391_ , \new_Sorter100|19392_ , \new_Sorter100|19393_ ,
    \new_Sorter100|19394_ , \new_Sorter100|19395_ , \new_Sorter100|19396_ ,
    \new_Sorter100|19397_ , \new_Sorter100|19398_ , \new_Sorter100|19400_ ,
    \new_Sorter100|19401_ , \new_Sorter100|19402_ , \new_Sorter100|19403_ ,
    \new_Sorter100|19404_ , \new_Sorter100|19405_ , \new_Sorter100|19406_ ,
    \new_Sorter100|19407_ , \new_Sorter100|19408_ , \new_Sorter100|19409_ ,
    \new_Sorter100|19410_ , \new_Sorter100|19411_ , \new_Sorter100|19412_ ,
    \new_Sorter100|19413_ , \new_Sorter100|19414_ , \new_Sorter100|19415_ ,
    \new_Sorter100|19416_ , \new_Sorter100|19417_ , \new_Sorter100|19418_ ,
    \new_Sorter100|19419_ , \new_Sorter100|19420_ , \new_Sorter100|19421_ ,
    \new_Sorter100|19422_ , \new_Sorter100|19423_ , \new_Sorter100|19424_ ,
    \new_Sorter100|19425_ , \new_Sorter100|19426_ , \new_Sorter100|19427_ ,
    \new_Sorter100|19428_ , \new_Sorter100|19429_ , \new_Sorter100|19430_ ,
    \new_Sorter100|19431_ , \new_Sorter100|19432_ , \new_Sorter100|19433_ ,
    \new_Sorter100|19434_ , \new_Sorter100|19435_ , \new_Sorter100|19436_ ,
    \new_Sorter100|19437_ , \new_Sorter100|19438_ , \new_Sorter100|19439_ ,
    \new_Sorter100|19440_ , \new_Sorter100|19441_ , \new_Sorter100|19442_ ,
    \new_Sorter100|19443_ , \new_Sorter100|19444_ , \new_Sorter100|19445_ ,
    \new_Sorter100|19446_ , \new_Sorter100|19447_ , \new_Sorter100|19448_ ,
    \new_Sorter100|19449_ , \new_Sorter100|19450_ , \new_Sorter100|19451_ ,
    \new_Sorter100|19452_ , \new_Sorter100|19453_ , \new_Sorter100|19454_ ,
    \new_Sorter100|19455_ , \new_Sorter100|19456_ , \new_Sorter100|19457_ ,
    \new_Sorter100|19458_ , \new_Sorter100|19459_ , \new_Sorter100|19460_ ,
    \new_Sorter100|19461_ , \new_Sorter100|19462_ , \new_Sorter100|19463_ ,
    \new_Sorter100|19464_ , \new_Sorter100|19465_ , \new_Sorter100|19466_ ,
    \new_Sorter100|19467_ , \new_Sorter100|19468_ , \new_Sorter100|19469_ ,
    \new_Sorter100|19470_ , \new_Sorter100|19471_ , \new_Sorter100|19472_ ,
    \new_Sorter100|19473_ , \new_Sorter100|19474_ , \new_Sorter100|19475_ ,
    \new_Sorter100|19476_ , \new_Sorter100|19477_ , \new_Sorter100|19478_ ,
    \new_Sorter100|19479_ , \new_Sorter100|19480_ , \new_Sorter100|19481_ ,
    \new_Sorter100|19482_ , \new_Sorter100|19483_ , \new_Sorter100|19484_ ,
    \new_Sorter100|19485_ , \new_Sorter100|19486_ , \new_Sorter100|19487_ ,
    \new_Sorter100|19488_ , \new_Sorter100|19489_ , \new_Sorter100|19490_ ,
    \new_Sorter100|19491_ , \new_Sorter100|19492_ , \new_Sorter100|19493_ ,
    \new_Sorter100|19494_ , \new_Sorter100|19495_ , \new_Sorter100|19496_ ,
    \new_Sorter100|19497_ , \new_Sorter100|19498_ , \new_Sorter100|19499_ ,
    \new_Sorter100|19500_ , \new_Sorter100|19599_ , \new_Sorter100|19501_ ,
    \new_Sorter100|19502_ , \new_Sorter100|19503_ , \new_Sorter100|19504_ ,
    \new_Sorter100|19505_ , \new_Sorter100|19506_ , \new_Sorter100|19507_ ,
    \new_Sorter100|19508_ , \new_Sorter100|19509_ , \new_Sorter100|19510_ ,
    \new_Sorter100|19511_ , \new_Sorter100|19512_ , \new_Sorter100|19513_ ,
    \new_Sorter100|19514_ , \new_Sorter100|19515_ , \new_Sorter100|19516_ ,
    \new_Sorter100|19517_ , \new_Sorter100|19518_ , \new_Sorter100|19519_ ,
    \new_Sorter100|19520_ , \new_Sorter100|19521_ , \new_Sorter100|19522_ ,
    \new_Sorter100|19523_ , \new_Sorter100|19524_ , \new_Sorter100|19525_ ,
    \new_Sorter100|19526_ , \new_Sorter100|19527_ , \new_Sorter100|19528_ ,
    \new_Sorter100|19529_ , \new_Sorter100|19530_ , \new_Sorter100|19531_ ,
    \new_Sorter100|19532_ , \new_Sorter100|19533_ , \new_Sorter100|19534_ ,
    \new_Sorter100|19535_ , \new_Sorter100|19536_ , \new_Sorter100|19537_ ,
    \new_Sorter100|19538_ , \new_Sorter100|19539_ , \new_Sorter100|19540_ ,
    \new_Sorter100|19541_ , \new_Sorter100|19542_ , \new_Sorter100|19543_ ,
    \new_Sorter100|19544_ , \new_Sorter100|19545_ , \new_Sorter100|19546_ ,
    \new_Sorter100|19547_ , \new_Sorter100|19548_ , \new_Sorter100|19549_ ,
    \new_Sorter100|19550_ , \new_Sorter100|19551_ , \new_Sorter100|19552_ ,
    \new_Sorter100|19553_ , \new_Sorter100|19554_ , \new_Sorter100|19555_ ,
    \new_Sorter100|19556_ , \new_Sorter100|19557_ , \new_Sorter100|19558_ ,
    \new_Sorter100|19559_ , \new_Sorter100|19560_ , \new_Sorter100|19561_ ,
    \new_Sorter100|19562_ , \new_Sorter100|19563_ , \new_Sorter100|19564_ ,
    \new_Sorter100|19565_ , \new_Sorter100|19566_ , \new_Sorter100|19567_ ,
    \new_Sorter100|19568_ , \new_Sorter100|19569_ , \new_Sorter100|19570_ ,
    \new_Sorter100|19571_ , \new_Sorter100|19572_ , \new_Sorter100|19573_ ,
    \new_Sorter100|19574_ , \new_Sorter100|19575_ , \new_Sorter100|19576_ ,
    \new_Sorter100|19577_ , \new_Sorter100|19578_ , \new_Sorter100|19579_ ,
    \new_Sorter100|19580_ , \new_Sorter100|19581_ , \new_Sorter100|19582_ ,
    \new_Sorter100|19583_ , \new_Sorter100|19584_ , \new_Sorter100|19585_ ,
    \new_Sorter100|19586_ , \new_Sorter100|19587_ , \new_Sorter100|19588_ ,
    \new_Sorter100|19589_ , \new_Sorter100|19590_ , \new_Sorter100|19591_ ,
    \new_Sorter100|19592_ , \new_Sorter100|19593_ , \new_Sorter100|19594_ ,
    \new_Sorter100|19595_ , \new_Sorter100|19596_ , \new_Sorter100|19597_ ,
    \new_Sorter100|19598_ , \new_Sorter100|19600_ , \new_Sorter100|19601_ ,
    \new_Sorter100|19602_ , \new_Sorter100|19603_ , \new_Sorter100|19604_ ,
    \new_Sorter100|19605_ , \new_Sorter100|19606_ , \new_Sorter100|19607_ ,
    \new_Sorter100|19608_ , \new_Sorter100|19609_ , \new_Sorter100|19610_ ,
    \new_Sorter100|19611_ , \new_Sorter100|19612_ , \new_Sorter100|19613_ ,
    \new_Sorter100|19614_ , \new_Sorter100|19615_ , \new_Sorter100|19616_ ,
    \new_Sorter100|19617_ , \new_Sorter100|19618_ , \new_Sorter100|19619_ ,
    \new_Sorter100|19620_ , \new_Sorter100|19621_ , \new_Sorter100|19622_ ,
    \new_Sorter100|19623_ , \new_Sorter100|19624_ , \new_Sorter100|19625_ ,
    \new_Sorter100|19626_ , \new_Sorter100|19627_ , \new_Sorter100|19628_ ,
    \new_Sorter100|19629_ , \new_Sorter100|19630_ , \new_Sorter100|19631_ ,
    \new_Sorter100|19632_ , \new_Sorter100|19633_ , \new_Sorter100|19634_ ,
    \new_Sorter100|19635_ , \new_Sorter100|19636_ , \new_Sorter100|19637_ ,
    \new_Sorter100|19638_ , \new_Sorter100|19639_ , \new_Sorter100|19640_ ,
    \new_Sorter100|19641_ , \new_Sorter100|19642_ , \new_Sorter100|19643_ ,
    \new_Sorter100|19644_ , \new_Sorter100|19645_ , \new_Sorter100|19646_ ,
    \new_Sorter100|19647_ , \new_Sorter100|19648_ , \new_Sorter100|19649_ ,
    \new_Sorter100|19650_ , \new_Sorter100|19651_ , \new_Sorter100|19652_ ,
    \new_Sorter100|19653_ , \new_Sorter100|19654_ , \new_Sorter100|19655_ ,
    \new_Sorter100|19656_ , \new_Sorter100|19657_ , \new_Sorter100|19658_ ,
    \new_Sorter100|19659_ , \new_Sorter100|19660_ , \new_Sorter100|19661_ ,
    \new_Sorter100|19662_ , \new_Sorter100|19663_ , \new_Sorter100|19664_ ,
    \new_Sorter100|19665_ , \new_Sorter100|19666_ , \new_Sorter100|19667_ ,
    \new_Sorter100|19668_ , \new_Sorter100|19669_ , \new_Sorter100|19670_ ,
    \new_Sorter100|19671_ , \new_Sorter100|19672_ , \new_Sorter100|19673_ ,
    \new_Sorter100|19674_ , \new_Sorter100|19675_ , \new_Sorter100|19676_ ,
    \new_Sorter100|19677_ , \new_Sorter100|19678_ , \new_Sorter100|19679_ ,
    \new_Sorter100|19680_ , \new_Sorter100|19681_ , \new_Sorter100|19682_ ,
    \new_Sorter100|19683_ , \new_Sorter100|19684_ , \new_Sorter100|19685_ ,
    \new_Sorter100|19686_ , \new_Sorter100|19687_ , \new_Sorter100|19688_ ,
    \new_Sorter100|19689_ , \new_Sorter100|19690_ , \new_Sorter100|19691_ ,
    \new_Sorter100|19692_ , \new_Sorter100|19693_ , \new_Sorter100|19694_ ,
    \new_Sorter100|19695_ , \new_Sorter100|19696_ , \new_Sorter100|19697_ ,
    \new_Sorter100|19698_ , \new_Sorter100|19699_ , \new_Sorter100|19700_ ,
    \new_Sorter100|19799_ , \new_Sorter100|19701_ , \new_Sorter100|19702_ ,
    \new_Sorter100|19703_ , \new_Sorter100|19704_ , \new_Sorter100|19705_ ,
    \new_Sorter100|19706_ , \new_Sorter100|19707_ , \new_Sorter100|19708_ ,
    \new_Sorter100|19709_ , \new_Sorter100|19710_ , \new_Sorter100|19711_ ,
    \new_Sorter100|19712_ , \new_Sorter100|19713_ , \new_Sorter100|19714_ ,
    \new_Sorter100|19715_ , \new_Sorter100|19716_ , \new_Sorter100|19717_ ,
    \new_Sorter100|19718_ , \new_Sorter100|19719_ , \new_Sorter100|19720_ ,
    \new_Sorter100|19721_ , \new_Sorter100|19722_ , \new_Sorter100|19723_ ,
    \new_Sorter100|19724_ , \new_Sorter100|19725_ , \new_Sorter100|19726_ ,
    \new_Sorter100|19727_ , \new_Sorter100|19728_ , \new_Sorter100|19729_ ,
    \new_Sorter100|19730_ , \new_Sorter100|19731_ , \new_Sorter100|19732_ ,
    \new_Sorter100|19733_ , \new_Sorter100|19734_ , \new_Sorter100|19735_ ,
    \new_Sorter100|19736_ , \new_Sorter100|19737_ , \new_Sorter100|19738_ ,
    \new_Sorter100|19739_ , \new_Sorter100|19740_ , \new_Sorter100|19741_ ,
    \new_Sorter100|19742_ , \new_Sorter100|19743_ , \new_Sorter100|19744_ ,
    \new_Sorter100|19745_ , \new_Sorter100|19746_ , \new_Sorter100|19747_ ,
    \new_Sorter100|19748_ , \new_Sorter100|19749_ , \new_Sorter100|19750_ ,
    \new_Sorter100|19751_ , \new_Sorter100|19752_ , \new_Sorter100|19753_ ,
    \new_Sorter100|19754_ , \new_Sorter100|19755_ , \new_Sorter100|19756_ ,
    \new_Sorter100|19757_ , \new_Sorter100|19758_ , \new_Sorter100|19759_ ,
    \new_Sorter100|19760_ , \new_Sorter100|19761_ , \new_Sorter100|19762_ ,
    \new_Sorter100|19763_ , \new_Sorter100|19764_ , \new_Sorter100|19765_ ,
    \new_Sorter100|19766_ , \new_Sorter100|19767_ , \new_Sorter100|19768_ ,
    \new_Sorter100|19769_ , \new_Sorter100|19770_ , \new_Sorter100|19771_ ,
    \new_Sorter100|19772_ , \new_Sorter100|19773_ , \new_Sorter100|19774_ ,
    \new_Sorter100|19775_ , \new_Sorter100|19776_ , \new_Sorter100|19777_ ,
    \new_Sorter100|19778_ , \new_Sorter100|19779_ , \new_Sorter100|19780_ ,
    \new_Sorter100|19781_ , \new_Sorter100|19782_ , \new_Sorter100|19783_ ,
    \new_Sorter100|19784_ , \new_Sorter100|19785_ , \new_Sorter100|19786_ ,
    \new_Sorter100|19787_ , \new_Sorter100|19788_ , \new_Sorter100|19789_ ,
    \new_Sorter100|19790_ , \new_Sorter100|19791_ , \new_Sorter100|19792_ ,
    \new_Sorter100|19793_ , \new_Sorter100|19794_ , \new_Sorter100|19795_ ,
    \new_Sorter100|19796_ , \new_Sorter100|19797_ , \new_Sorter100|19798_ ;
  assign \new_Sorter100|0000_  = x00 & x01;
  assign \new_Sorter100|0001_  = x00 | x01;
  assign \new_Sorter100|0002_  = x02 & x03;
  assign \new_Sorter100|0003_  = x02 | x03;
  assign \new_Sorter100|0004_  = x04 & x05;
  assign \new_Sorter100|0005_  = x04 | x05;
  assign \new_Sorter100|0006_  = x06 & x07;
  assign \new_Sorter100|0007_  = x06 | x07;
  assign \new_Sorter100|0008_  = x08 & x09;
  assign \new_Sorter100|0009_  = x08 | x09;
  assign \new_Sorter100|0010_  = x10 & x11;
  assign \new_Sorter100|0011_  = x10 | x11;
  assign \new_Sorter100|0012_  = x12 & x13;
  assign \new_Sorter100|0013_  = x12 | x13;
  assign \new_Sorter100|0014_  = x14 & x15;
  assign \new_Sorter100|0015_  = x14 | x15;
  assign \new_Sorter100|0016_  = x16 & x17;
  assign \new_Sorter100|0017_  = x16 | x17;
  assign \new_Sorter100|0018_  = x18 & x19;
  assign \new_Sorter100|0019_  = x18 | x19;
  assign \new_Sorter100|0020_  = x20 & x21;
  assign \new_Sorter100|0021_  = x20 | x21;
  assign \new_Sorter100|0022_  = x22 & x23;
  assign \new_Sorter100|0023_  = x22 | x23;
  assign \new_Sorter100|0024_  = x24 & x25;
  assign \new_Sorter100|0025_  = x24 | x25;
  assign \new_Sorter100|0026_  = x26 & x27;
  assign \new_Sorter100|0027_  = x26 | x27;
  assign \new_Sorter100|0028_  = x28 & x29;
  assign \new_Sorter100|0029_  = x28 | x29;
  assign \new_Sorter100|0030_  = x30 & x31;
  assign \new_Sorter100|0031_  = x30 | x31;
  assign \new_Sorter100|0032_  = x32 & x33;
  assign \new_Sorter100|0033_  = x32 | x33;
  assign \new_Sorter100|0034_  = x34 & x35;
  assign \new_Sorter100|0035_  = x34 | x35;
  assign \new_Sorter100|0036_  = x36 & x37;
  assign \new_Sorter100|0037_  = x36 | x37;
  assign \new_Sorter100|0038_  = x38 & x39;
  assign \new_Sorter100|0039_  = x38 | x39;
  assign \new_Sorter100|0040_  = x40 & x41;
  assign \new_Sorter100|0041_  = x40 | x41;
  assign \new_Sorter100|0042_  = x42 & x43;
  assign \new_Sorter100|0043_  = x42 | x43;
  assign \new_Sorter100|0044_  = x44 & x45;
  assign \new_Sorter100|0045_  = x44 | x45;
  assign \new_Sorter100|0046_  = x46 & x47;
  assign \new_Sorter100|0047_  = x46 | x47;
  assign \new_Sorter100|0048_  = x48 & x49;
  assign \new_Sorter100|0049_  = x48 | x49;
  assign \new_Sorter100|0050_  = x50 & x51;
  assign \new_Sorter100|0051_  = x50 | x51;
  assign \new_Sorter100|0052_  = x52 & x53;
  assign \new_Sorter100|0053_  = x52 | x53;
  assign \new_Sorter100|0054_  = x54 & x55;
  assign \new_Sorter100|0055_  = x54 | x55;
  assign \new_Sorter100|0056_  = x56 & x57;
  assign \new_Sorter100|0057_  = x56 | x57;
  assign \new_Sorter100|0058_  = x58 & x59;
  assign \new_Sorter100|0059_  = x58 | x59;
  assign \new_Sorter100|0060_  = x60 & x61;
  assign \new_Sorter100|0061_  = x60 | x61;
  assign \new_Sorter100|0062_  = x62 & x63;
  assign \new_Sorter100|0063_  = x62 | x63;
  assign \new_Sorter100|0064_  = x64 & x65;
  assign \new_Sorter100|0065_  = x64 | x65;
  assign \new_Sorter100|0066_  = x66 & x67;
  assign \new_Sorter100|0067_  = x66 | x67;
  assign \new_Sorter100|0068_  = x68 & x69;
  assign \new_Sorter100|0069_  = x68 | x69;
  assign \new_Sorter100|0070_  = x70 & x71;
  assign \new_Sorter100|0071_  = x70 | x71;
  assign \new_Sorter100|0072_  = x72 & x73;
  assign \new_Sorter100|0073_  = x72 | x73;
  assign \new_Sorter100|0074_  = x74 & x75;
  assign \new_Sorter100|0075_  = x74 | x75;
  assign \new_Sorter100|0076_  = x76 & x77;
  assign \new_Sorter100|0077_  = x76 | x77;
  assign \new_Sorter100|0078_  = x78 & x79;
  assign \new_Sorter100|0079_  = x78 | x79;
  assign \new_Sorter100|0080_  = x80 & x81;
  assign \new_Sorter100|0081_  = x80 | x81;
  assign \new_Sorter100|0082_  = x82 & x83;
  assign \new_Sorter100|0083_  = x82 | x83;
  assign \new_Sorter100|0084_  = x84 & x85;
  assign \new_Sorter100|0085_  = x84 | x85;
  assign \new_Sorter100|0086_  = x86 & x87;
  assign \new_Sorter100|0087_  = x86 | x87;
  assign \new_Sorter100|0088_  = x88 & x89;
  assign \new_Sorter100|0089_  = x88 | x89;
  assign \new_Sorter100|0090_  = x90 & x91;
  assign \new_Sorter100|0091_  = x90 | x91;
  assign \new_Sorter100|0092_  = x92 & x93;
  assign \new_Sorter100|0093_  = x92 | x93;
  assign \new_Sorter100|0094_  = x94 & x95;
  assign \new_Sorter100|0095_  = x94 | x95;
  assign \new_Sorter100|0096_  = x96 & x97;
  assign \new_Sorter100|0097_  = x96 | x97;
  assign \new_Sorter100|0098_  = x98 & x99;
  assign \new_Sorter100|0099_  = x98 | x99;
  assign \new_Sorter100|0100_  = \new_Sorter100|0000_ ;
  assign \new_Sorter100|0199_  = \new_Sorter100|0099_ ;
  assign \new_Sorter100|0101_  = \new_Sorter100|0001_  & \new_Sorter100|0002_ ;
  assign \new_Sorter100|0102_  = \new_Sorter100|0001_  | \new_Sorter100|0002_ ;
  assign \new_Sorter100|0103_  = \new_Sorter100|0003_  & \new_Sorter100|0004_ ;
  assign \new_Sorter100|0104_  = \new_Sorter100|0003_  | \new_Sorter100|0004_ ;
  assign \new_Sorter100|0105_  = \new_Sorter100|0005_  & \new_Sorter100|0006_ ;
  assign \new_Sorter100|0106_  = \new_Sorter100|0005_  | \new_Sorter100|0006_ ;
  assign \new_Sorter100|0107_  = \new_Sorter100|0007_  & \new_Sorter100|0008_ ;
  assign \new_Sorter100|0108_  = \new_Sorter100|0007_  | \new_Sorter100|0008_ ;
  assign \new_Sorter100|0109_  = \new_Sorter100|0009_  & \new_Sorter100|0010_ ;
  assign \new_Sorter100|0110_  = \new_Sorter100|0009_  | \new_Sorter100|0010_ ;
  assign \new_Sorter100|0111_  = \new_Sorter100|0011_  & \new_Sorter100|0012_ ;
  assign \new_Sorter100|0112_  = \new_Sorter100|0011_  | \new_Sorter100|0012_ ;
  assign \new_Sorter100|0113_  = \new_Sorter100|0013_  & \new_Sorter100|0014_ ;
  assign \new_Sorter100|0114_  = \new_Sorter100|0013_  | \new_Sorter100|0014_ ;
  assign \new_Sorter100|0115_  = \new_Sorter100|0015_  & \new_Sorter100|0016_ ;
  assign \new_Sorter100|0116_  = \new_Sorter100|0015_  | \new_Sorter100|0016_ ;
  assign \new_Sorter100|0117_  = \new_Sorter100|0017_  & \new_Sorter100|0018_ ;
  assign \new_Sorter100|0118_  = \new_Sorter100|0017_  | \new_Sorter100|0018_ ;
  assign \new_Sorter100|0119_  = \new_Sorter100|0019_  & \new_Sorter100|0020_ ;
  assign \new_Sorter100|0120_  = \new_Sorter100|0019_  | \new_Sorter100|0020_ ;
  assign \new_Sorter100|0121_  = \new_Sorter100|0021_  & \new_Sorter100|0022_ ;
  assign \new_Sorter100|0122_  = \new_Sorter100|0021_  | \new_Sorter100|0022_ ;
  assign \new_Sorter100|0123_  = \new_Sorter100|0023_  & \new_Sorter100|0024_ ;
  assign \new_Sorter100|0124_  = \new_Sorter100|0023_  | \new_Sorter100|0024_ ;
  assign \new_Sorter100|0125_  = \new_Sorter100|0025_  & \new_Sorter100|0026_ ;
  assign \new_Sorter100|0126_  = \new_Sorter100|0025_  | \new_Sorter100|0026_ ;
  assign \new_Sorter100|0127_  = \new_Sorter100|0027_  & \new_Sorter100|0028_ ;
  assign \new_Sorter100|0128_  = \new_Sorter100|0027_  | \new_Sorter100|0028_ ;
  assign \new_Sorter100|0129_  = \new_Sorter100|0029_  & \new_Sorter100|0030_ ;
  assign \new_Sorter100|0130_  = \new_Sorter100|0029_  | \new_Sorter100|0030_ ;
  assign \new_Sorter100|0131_  = \new_Sorter100|0031_  & \new_Sorter100|0032_ ;
  assign \new_Sorter100|0132_  = \new_Sorter100|0031_  | \new_Sorter100|0032_ ;
  assign \new_Sorter100|0133_  = \new_Sorter100|0033_  & \new_Sorter100|0034_ ;
  assign \new_Sorter100|0134_  = \new_Sorter100|0033_  | \new_Sorter100|0034_ ;
  assign \new_Sorter100|0135_  = \new_Sorter100|0035_  & \new_Sorter100|0036_ ;
  assign \new_Sorter100|0136_  = \new_Sorter100|0035_  | \new_Sorter100|0036_ ;
  assign \new_Sorter100|0137_  = \new_Sorter100|0037_  & \new_Sorter100|0038_ ;
  assign \new_Sorter100|0138_  = \new_Sorter100|0037_  | \new_Sorter100|0038_ ;
  assign \new_Sorter100|0139_  = \new_Sorter100|0039_  & \new_Sorter100|0040_ ;
  assign \new_Sorter100|0140_  = \new_Sorter100|0039_  | \new_Sorter100|0040_ ;
  assign \new_Sorter100|0141_  = \new_Sorter100|0041_  & \new_Sorter100|0042_ ;
  assign \new_Sorter100|0142_  = \new_Sorter100|0041_  | \new_Sorter100|0042_ ;
  assign \new_Sorter100|0143_  = \new_Sorter100|0043_  & \new_Sorter100|0044_ ;
  assign \new_Sorter100|0144_  = \new_Sorter100|0043_  | \new_Sorter100|0044_ ;
  assign \new_Sorter100|0145_  = \new_Sorter100|0045_  & \new_Sorter100|0046_ ;
  assign \new_Sorter100|0146_  = \new_Sorter100|0045_  | \new_Sorter100|0046_ ;
  assign \new_Sorter100|0147_  = \new_Sorter100|0047_  & \new_Sorter100|0048_ ;
  assign \new_Sorter100|0148_  = \new_Sorter100|0047_  | \new_Sorter100|0048_ ;
  assign \new_Sorter100|0149_  = \new_Sorter100|0049_  & \new_Sorter100|0050_ ;
  assign \new_Sorter100|0150_  = \new_Sorter100|0049_  | \new_Sorter100|0050_ ;
  assign \new_Sorter100|0151_  = \new_Sorter100|0051_  & \new_Sorter100|0052_ ;
  assign \new_Sorter100|0152_  = \new_Sorter100|0051_  | \new_Sorter100|0052_ ;
  assign \new_Sorter100|0153_  = \new_Sorter100|0053_  & \new_Sorter100|0054_ ;
  assign \new_Sorter100|0154_  = \new_Sorter100|0053_  | \new_Sorter100|0054_ ;
  assign \new_Sorter100|0155_  = \new_Sorter100|0055_  & \new_Sorter100|0056_ ;
  assign \new_Sorter100|0156_  = \new_Sorter100|0055_  | \new_Sorter100|0056_ ;
  assign \new_Sorter100|0157_  = \new_Sorter100|0057_  & \new_Sorter100|0058_ ;
  assign \new_Sorter100|0158_  = \new_Sorter100|0057_  | \new_Sorter100|0058_ ;
  assign \new_Sorter100|0159_  = \new_Sorter100|0059_  & \new_Sorter100|0060_ ;
  assign \new_Sorter100|0160_  = \new_Sorter100|0059_  | \new_Sorter100|0060_ ;
  assign \new_Sorter100|0161_  = \new_Sorter100|0061_  & \new_Sorter100|0062_ ;
  assign \new_Sorter100|0162_  = \new_Sorter100|0061_  | \new_Sorter100|0062_ ;
  assign \new_Sorter100|0163_  = \new_Sorter100|0063_  & \new_Sorter100|0064_ ;
  assign \new_Sorter100|0164_  = \new_Sorter100|0063_  | \new_Sorter100|0064_ ;
  assign \new_Sorter100|0165_  = \new_Sorter100|0065_  & \new_Sorter100|0066_ ;
  assign \new_Sorter100|0166_  = \new_Sorter100|0065_  | \new_Sorter100|0066_ ;
  assign \new_Sorter100|0167_  = \new_Sorter100|0067_  & \new_Sorter100|0068_ ;
  assign \new_Sorter100|0168_  = \new_Sorter100|0067_  | \new_Sorter100|0068_ ;
  assign \new_Sorter100|0169_  = \new_Sorter100|0069_  & \new_Sorter100|0070_ ;
  assign \new_Sorter100|0170_  = \new_Sorter100|0069_  | \new_Sorter100|0070_ ;
  assign \new_Sorter100|0171_  = \new_Sorter100|0071_  & \new_Sorter100|0072_ ;
  assign \new_Sorter100|0172_  = \new_Sorter100|0071_  | \new_Sorter100|0072_ ;
  assign \new_Sorter100|0173_  = \new_Sorter100|0073_  & \new_Sorter100|0074_ ;
  assign \new_Sorter100|0174_  = \new_Sorter100|0073_  | \new_Sorter100|0074_ ;
  assign \new_Sorter100|0175_  = \new_Sorter100|0075_  & \new_Sorter100|0076_ ;
  assign \new_Sorter100|0176_  = \new_Sorter100|0075_  | \new_Sorter100|0076_ ;
  assign \new_Sorter100|0177_  = \new_Sorter100|0077_  & \new_Sorter100|0078_ ;
  assign \new_Sorter100|0178_  = \new_Sorter100|0077_  | \new_Sorter100|0078_ ;
  assign \new_Sorter100|0179_  = \new_Sorter100|0079_  & \new_Sorter100|0080_ ;
  assign \new_Sorter100|0180_  = \new_Sorter100|0079_  | \new_Sorter100|0080_ ;
  assign \new_Sorter100|0181_  = \new_Sorter100|0081_  & \new_Sorter100|0082_ ;
  assign \new_Sorter100|0182_  = \new_Sorter100|0081_  | \new_Sorter100|0082_ ;
  assign \new_Sorter100|0183_  = \new_Sorter100|0083_  & \new_Sorter100|0084_ ;
  assign \new_Sorter100|0184_  = \new_Sorter100|0083_  | \new_Sorter100|0084_ ;
  assign \new_Sorter100|0185_  = \new_Sorter100|0085_  & \new_Sorter100|0086_ ;
  assign \new_Sorter100|0186_  = \new_Sorter100|0085_  | \new_Sorter100|0086_ ;
  assign \new_Sorter100|0187_  = \new_Sorter100|0087_  & \new_Sorter100|0088_ ;
  assign \new_Sorter100|0188_  = \new_Sorter100|0087_  | \new_Sorter100|0088_ ;
  assign \new_Sorter100|0189_  = \new_Sorter100|0089_  & \new_Sorter100|0090_ ;
  assign \new_Sorter100|0190_  = \new_Sorter100|0089_  | \new_Sorter100|0090_ ;
  assign \new_Sorter100|0191_  = \new_Sorter100|0091_  & \new_Sorter100|0092_ ;
  assign \new_Sorter100|0192_  = \new_Sorter100|0091_  | \new_Sorter100|0092_ ;
  assign \new_Sorter100|0193_  = \new_Sorter100|0093_  & \new_Sorter100|0094_ ;
  assign \new_Sorter100|0194_  = \new_Sorter100|0093_  | \new_Sorter100|0094_ ;
  assign \new_Sorter100|0195_  = \new_Sorter100|0095_  & \new_Sorter100|0096_ ;
  assign \new_Sorter100|0196_  = \new_Sorter100|0095_  | \new_Sorter100|0096_ ;
  assign \new_Sorter100|0197_  = \new_Sorter100|0097_  & \new_Sorter100|0098_ ;
  assign \new_Sorter100|0198_  = \new_Sorter100|0097_  | \new_Sorter100|0098_ ;
  assign \new_Sorter100|0200_  = \new_Sorter100|0100_  & \new_Sorter100|0101_ ;
  assign \new_Sorter100|0201_  = \new_Sorter100|0100_  | \new_Sorter100|0101_ ;
  assign \new_Sorter100|0202_  = \new_Sorter100|0102_  & \new_Sorter100|0103_ ;
  assign \new_Sorter100|0203_  = \new_Sorter100|0102_  | \new_Sorter100|0103_ ;
  assign \new_Sorter100|0204_  = \new_Sorter100|0104_  & \new_Sorter100|0105_ ;
  assign \new_Sorter100|0205_  = \new_Sorter100|0104_  | \new_Sorter100|0105_ ;
  assign \new_Sorter100|0206_  = \new_Sorter100|0106_  & \new_Sorter100|0107_ ;
  assign \new_Sorter100|0207_  = \new_Sorter100|0106_  | \new_Sorter100|0107_ ;
  assign \new_Sorter100|0208_  = \new_Sorter100|0108_  & \new_Sorter100|0109_ ;
  assign \new_Sorter100|0209_  = \new_Sorter100|0108_  | \new_Sorter100|0109_ ;
  assign \new_Sorter100|0210_  = \new_Sorter100|0110_  & \new_Sorter100|0111_ ;
  assign \new_Sorter100|0211_  = \new_Sorter100|0110_  | \new_Sorter100|0111_ ;
  assign \new_Sorter100|0212_  = \new_Sorter100|0112_  & \new_Sorter100|0113_ ;
  assign \new_Sorter100|0213_  = \new_Sorter100|0112_  | \new_Sorter100|0113_ ;
  assign \new_Sorter100|0214_  = \new_Sorter100|0114_  & \new_Sorter100|0115_ ;
  assign \new_Sorter100|0215_  = \new_Sorter100|0114_  | \new_Sorter100|0115_ ;
  assign \new_Sorter100|0216_  = \new_Sorter100|0116_  & \new_Sorter100|0117_ ;
  assign \new_Sorter100|0217_  = \new_Sorter100|0116_  | \new_Sorter100|0117_ ;
  assign \new_Sorter100|0218_  = \new_Sorter100|0118_  & \new_Sorter100|0119_ ;
  assign \new_Sorter100|0219_  = \new_Sorter100|0118_  | \new_Sorter100|0119_ ;
  assign \new_Sorter100|0220_  = \new_Sorter100|0120_  & \new_Sorter100|0121_ ;
  assign \new_Sorter100|0221_  = \new_Sorter100|0120_  | \new_Sorter100|0121_ ;
  assign \new_Sorter100|0222_  = \new_Sorter100|0122_  & \new_Sorter100|0123_ ;
  assign \new_Sorter100|0223_  = \new_Sorter100|0122_  | \new_Sorter100|0123_ ;
  assign \new_Sorter100|0224_  = \new_Sorter100|0124_  & \new_Sorter100|0125_ ;
  assign \new_Sorter100|0225_  = \new_Sorter100|0124_  | \new_Sorter100|0125_ ;
  assign \new_Sorter100|0226_  = \new_Sorter100|0126_  & \new_Sorter100|0127_ ;
  assign \new_Sorter100|0227_  = \new_Sorter100|0126_  | \new_Sorter100|0127_ ;
  assign \new_Sorter100|0228_  = \new_Sorter100|0128_  & \new_Sorter100|0129_ ;
  assign \new_Sorter100|0229_  = \new_Sorter100|0128_  | \new_Sorter100|0129_ ;
  assign \new_Sorter100|0230_  = \new_Sorter100|0130_  & \new_Sorter100|0131_ ;
  assign \new_Sorter100|0231_  = \new_Sorter100|0130_  | \new_Sorter100|0131_ ;
  assign \new_Sorter100|0232_  = \new_Sorter100|0132_  & \new_Sorter100|0133_ ;
  assign \new_Sorter100|0233_  = \new_Sorter100|0132_  | \new_Sorter100|0133_ ;
  assign \new_Sorter100|0234_  = \new_Sorter100|0134_  & \new_Sorter100|0135_ ;
  assign \new_Sorter100|0235_  = \new_Sorter100|0134_  | \new_Sorter100|0135_ ;
  assign \new_Sorter100|0236_  = \new_Sorter100|0136_  & \new_Sorter100|0137_ ;
  assign \new_Sorter100|0237_  = \new_Sorter100|0136_  | \new_Sorter100|0137_ ;
  assign \new_Sorter100|0238_  = \new_Sorter100|0138_  & \new_Sorter100|0139_ ;
  assign \new_Sorter100|0239_  = \new_Sorter100|0138_  | \new_Sorter100|0139_ ;
  assign \new_Sorter100|0240_  = \new_Sorter100|0140_  & \new_Sorter100|0141_ ;
  assign \new_Sorter100|0241_  = \new_Sorter100|0140_  | \new_Sorter100|0141_ ;
  assign \new_Sorter100|0242_  = \new_Sorter100|0142_  & \new_Sorter100|0143_ ;
  assign \new_Sorter100|0243_  = \new_Sorter100|0142_  | \new_Sorter100|0143_ ;
  assign \new_Sorter100|0244_  = \new_Sorter100|0144_  & \new_Sorter100|0145_ ;
  assign \new_Sorter100|0245_  = \new_Sorter100|0144_  | \new_Sorter100|0145_ ;
  assign \new_Sorter100|0246_  = \new_Sorter100|0146_  & \new_Sorter100|0147_ ;
  assign \new_Sorter100|0247_  = \new_Sorter100|0146_  | \new_Sorter100|0147_ ;
  assign \new_Sorter100|0248_  = \new_Sorter100|0148_  & \new_Sorter100|0149_ ;
  assign \new_Sorter100|0249_  = \new_Sorter100|0148_  | \new_Sorter100|0149_ ;
  assign \new_Sorter100|0250_  = \new_Sorter100|0150_  & \new_Sorter100|0151_ ;
  assign \new_Sorter100|0251_  = \new_Sorter100|0150_  | \new_Sorter100|0151_ ;
  assign \new_Sorter100|0252_  = \new_Sorter100|0152_  & \new_Sorter100|0153_ ;
  assign \new_Sorter100|0253_  = \new_Sorter100|0152_  | \new_Sorter100|0153_ ;
  assign \new_Sorter100|0254_  = \new_Sorter100|0154_  & \new_Sorter100|0155_ ;
  assign \new_Sorter100|0255_  = \new_Sorter100|0154_  | \new_Sorter100|0155_ ;
  assign \new_Sorter100|0256_  = \new_Sorter100|0156_  & \new_Sorter100|0157_ ;
  assign \new_Sorter100|0257_  = \new_Sorter100|0156_  | \new_Sorter100|0157_ ;
  assign \new_Sorter100|0258_  = \new_Sorter100|0158_  & \new_Sorter100|0159_ ;
  assign \new_Sorter100|0259_  = \new_Sorter100|0158_  | \new_Sorter100|0159_ ;
  assign \new_Sorter100|0260_  = \new_Sorter100|0160_  & \new_Sorter100|0161_ ;
  assign \new_Sorter100|0261_  = \new_Sorter100|0160_  | \new_Sorter100|0161_ ;
  assign \new_Sorter100|0262_  = \new_Sorter100|0162_  & \new_Sorter100|0163_ ;
  assign \new_Sorter100|0263_  = \new_Sorter100|0162_  | \new_Sorter100|0163_ ;
  assign \new_Sorter100|0264_  = \new_Sorter100|0164_  & \new_Sorter100|0165_ ;
  assign \new_Sorter100|0265_  = \new_Sorter100|0164_  | \new_Sorter100|0165_ ;
  assign \new_Sorter100|0266_  = \new_Sorter100|0166_  & \new_Sorter100|0167_ ;
  assign \new_Sorter100|0267_  = \new_Sorter100|0166_  | \new_Sorter100|0167_ ;
  assign \new_Sorter100|0268_  = \new_Sorter100|0168_  & \new_Sorter100|0169_ ;
  assign \new_Sorter100|0269_  = \new_Sorter100|0168_  | \new_Sorter100|0169_ ;
  assign \new_Sorter100|0270_  = \new_Sorter100|0170_  & \new_Sorter100|0171_ ;
  assign \new_Sorter100|0271_  = \new_Sorter100|0170_  | \new_Sorter100|0171_ ;
  assign \new_Sorter100|0272_  = \new_Sorter100|0172_  & \new_Sorter100|0173_ ;
  assign \new_Sorter100|0273_  = \new_Sorter100|0172_  | \new_Sorter100|0173_ ;
  assign \new_Sorter100|0274_  = \new_Sorter100|0174_  & \new_Sorter100|0175_ ;
  assign \new_Sorter100|0275_  = \new_Sorter100|0174_  | \new_Sorter100|0175_ ;
  assign \new_Sorter100|0276_  = \new_Sorter100|0176_  & \new_Sorter100|0177_ ;
  assign \new_Sorter100|0277_  = \new_Sorter100|0176_  | \new_Sorter100|0177_ ;
  assign \new_Sorter100|0278_  = \new_Sorter100|0178_  & \new_Sorter100|0179_ ;
  assign \new_Sorter100|0279_  = \new_Sorter100|0178_  | \new_Sorter100|0179_ ;
  assign \new_Sorter100|0280_  = \new_Sorter100|0180_  & \new_Sorter100|0181_ ;
  assign \new_Sorter100|0281_  = \new_Sorter100|0180_  | \new_Sorter100|0181_ ;
  assign \new_Sorter100|0282_  = \new_Sorter100|0182_  & \new_Sorter100|0183_ ;
  assign \new_Sorter100|0283_  = \new_Sorter100|0182_  | \new_Sorter100|0183_ ;
  assign \new_Sorter100|0284_  = \new_Sorter100|0184_  & \new_Sorter100|0185_ ;
  assign \new_Sorter100|0285_  = \new_Sorter100|0184_  | \new_Sorter100|0185_ ;
  assign \new_Sorter100|0286_  = \new_Sorter100|0186_  & \new_Sorter100|0187_ ;
  assign \new_Sorter100|0287_  = \new_Sorter100|0186_  | \new_Sorter100|0187_ ;
  assign \new_Sorter100|0288_  = \new_Sorter100|0188_  & \new_Sorter100|0189_ ;
  assign \new_Sorter100|0289_  = \new_Sorter100|0188_  | \new_Sorter100|0189_ ;
  assign \new_Sorter100|0290_  = \new_Sorter100|0190_  & \new_Sorter100|0191_ ;
  assign \new_Sorter100|0291_  = \new_Sorter100|0190_  | \new_Sorter100|0191_ ;
  assign \new_Sorter100|0292_  = \new_Sorter100|0192_  & \new_Sorter100|0193_ ;
  assign \new_Sorter100|0293_  = \new_Sorter100|0192_  | \new_Sorter100|0193_ ;
  assign \new_Sorter100|0294_  = \new_Sorter100|0194_  & \new_Sorter100|0195_ ;
  assign \new_Sorter100|0295_  = \new_Sorter100|0194_  | \new_Sorter100|0195_ ;
  assign \new_Sorter100|0296_  = \new_Sorter100|0196_  & \new_Sorter100|0197_ ;
  assign \new_Sorter100|0297_  = \new_Sorter100|0196_  | \new_Sorter100|0197_ ;
  assign \new_Sorter100|0298_  = \new_Sorter100|0198_  & \new_Sorter100|0199_ ;
  assign \new_Sorter100|0299_  = \new_Sorter100|0198_  | \new_Sorter100|0199_ ;
  assign \new_Sorter100|0300_  = \new_Sorter100|0200_ ;
  assign \new_Sorter100|0399_  = \new_Sorter100|0299_ ;
  assign \new_Sorter100|0301_  = \new_Sorter100|0201_  & \new_Sorter100|0202_ ;
  assign \new_Sorter100|0302_  = \new_Sorter100|0201_  | \new_Sorter100|0202_ ;
  assign \new_Sorter100|0303_  = \new_Sorter100|0203_  & \new_Sorter100|0204_ ;
  assign \new_Sorter100|0304_  = \new_Sorter100|0203_  | \new_Sorter100|0204_ ;
  assign \new_Sorter100|0305_  = \new_Sorter100|0205_  & \new_Sorter100|0206_ ;
  assign \new_Sorter100|0306_  = \new_Sorter100|0205_  | \new_Sorter100|0206_ ;
  assign \new_Sorter100|0307_  = \new_Sorter100|0207_  & \new_Sorter100|0208_ ;
  assign \new_Sorter100|0308_  = \new_Sorter100|0207_  | \new_Sorter100|0208_ ;
  assign \new_Sorter100|0309_  = \new_Sorter100|0209_  & \new_Sorter100|0210_ ;
  assign \new_Sorter100|0310_  = \new_Sorter100|0209_  | \new_Sorter100|0210_ ;
  assign \new_Sorter100|0311_  = \new_Sorter100|0211_  & \new_Sorter100|0212_ ;
  assign \new_Sorter100|0312_  = \new_Sorter100|0211_  | \new_Sorter100|0212_ ;
  assign \new_Sorter100|0313_  = \new_Sorter100|0213_  & \new_Sorter100|0214_ ;
  assign \new_Sorter100|0314_  = \new_Sorter100|0213_  | \new_Sorter100|0214_ ;
  assign \new_Sorter100|0315_  = \new_Sorter100|0215_  & \new_Sorter100|0216_ ;
  assign \new_Sorter100|0316_  = \new_Sorter100|0215_  | \new_Sorter100|0216_ ;
  assign \new_Sorter100|0317_  = \new_Sorter100|0217_  & \new_Sorter100|0218_ ;
  assign \new_Sorter100|0318_  = \new_Sorter100|0217_  | \new_Sorter100|0218_ ;
  assign \new_Sorter100|0319_  = \new_Sorter100|0219_  & \new_Sorter100|0220_ ;
  assign \new_Sorter100|0320_  = \new_Sorter100|0219_  | \new_Sorter100|0220_ ;
  assign \new_Sorter100|0321_  = \new_Sorter100|0221_  & \new_Sorter100|0222_ ;
  assign \new_Sorter100|0322_  = \new_Sorter100|0221_  | \new_Sorter100|0222_ ;
  assign \new_Sorter100|0323_  = \new_Sorter100|0223_  & \new_Sorter100|0224_ ;
  assign \new_Sorter100|0324_  = \new_Sorter100|0223_  | \new_Sorter100|0224_ ;
  assign \new_Sorter100|0325_  = \new_Sorter100|0225_  & \new_Sorter100|0226_ ;
  assign \new_Sorter100|0326_  = \new_Sorter100|0225_  | \new_Sorter100|0226_ ;
  assign \new_Sorter100|0327_  = \new_Sorter100|0227_  & \new_Sorter100|0228_ ;
  assign \new_Sorter100|0328_  = \new_Sorter100|0227_  | \new_Sorter100|0228_ ;
  assign \new_Sorter100|0329_  = \new_Sorter100|0229_  & \new_Sorter100|0230_ ;
  assign \new_Sorter100|0330_  = \new_Sorter100|0229_  | \new_Sorter100|0230_ ;
  assign \new_Sorter100|0331_  = \new_Sorter100|0231_  & \new_Sorter100|0232_ ;
  assign \new_Sorter100|0332_  = \new_Sorter100|0231_  | \new_Sorter100|0232_ ;
  assign \new_Sorter100|0333_  = \new_Sorter100|0233_  & \new_Sorter100|0234_ ;
  assign \new_Sorter100|0334_  = \new_Sorter100|0233_  | \new_Sorter100|0234_ ;
  assign \new_Sorter100|0335_  = \new_Sorter100|0235_  & \new_Sorter100|0236_ ;
  assign \new_Sorter100|0336_  = \new_Sorter100|0235_  | \new_Sorter100|0236_ ;
  assign \new_Sorter100|0337_  = \new_Sorter100|0237_  & \new_Sorter100|0238_ ;
  assign \new_Sorter100|0338_  = \new_Sorter100|0237_  | \new_Sorter100|0238_ ;
  assign \new_Sorter100|0339_  = \new_Sorter100|0239_  & \new_Sorter100|0240_ ;
  assign \new_Sorter100|0340_  = \new_Sorter100|0239_  | \new_Sorter100|0240_ ;
  assign \new_Sorter100|0341_  = \new_Sorter100|0241_  & \new_Sorter100|0242_ ;
  assign \new_Sorter100|0342_  = \new_Sorter100|0241_  | \new_Sorter100|0242_ ;
  assign \new_Sorter100|0343_  = \new_Sorter100|0243_  & \new_Sorter100|0244_ ;
  assign \new_Sorter100|0344_  = \new_Sorter100|0243_  | \new_Sorter100|0244_ ;
  assign \new_Sorter100|0345_  = \new_Sorter100|0245_  & \new_Sorter100|0246_ ;
  assign \new_Sorter100|0346_  = \new_Sorter100|0245_  | \new_Sorter100|0246_ ;
  assign \new_Sorter100|0347_  = \new_Sorter100|0247_  & \new_Sorter100|0248_ ;
  assign \new_Sorter100|0348_  = \new_Sorter100|0247_  | \new_Sorter100|0248_ ;
  assign \new_Sorter100|0349_  = \new_Sorter100|0249_  & \new_Sorter100|0250_ ;
  assign \new_Sorter100|0350_  = \new_Sorter100|0249_  | \new_Sorter100|0250_ ;
  assign \new_Sorter100|0351_  = \new_Sorter100|0251_  & \new_Sorter100|0252_ ;
  assign \new_Sorter100|0352_  = \new_Sorter100|0251_  | \new_Sorter100|0252_ ;
  assign \new_Sorter100|0353_  = \new_Sorter100|0253_  & \new_Sorter100|0254_ ;
  assign \new_Sorter100|0354_  = \new_Sorter100|0253_  | \new_Sorter100|0254_ ;
  assign \new_Sorter100|0355_  = \new_Sorter100|0255_  & \new_Sorter100|0256_ ;
  assign \new_Sorter100|0356_  = \new_Sorter100|0255_  | \new_Sorter100|0256_ ;
  assign \new_Sorter100|0357_  = \new_Sorter100|0257_  & \new_Sorter100|0258_ ;
  assign \new_Sorter100|0358_  = \new_Sorter100|0257_  | \new_Sorter100|0258_ ;
  assign \new_Sorter100|0359_  = \new_Sorter100|0259_  & \new_Sorter100|0260_ ;
  assign \new_Sorter100|0360_  = \new_Sorter100|0259_  | \new_Sorter100|0260_ ;
  assign \new_Sorter100|0361_  = \new_Sorter100|0261_  & \new_Sorter100|0262_ ;
  assign \new_Sorter100|0362_  = \new_Sorter100|0261_  | \new_Sorter100|0262_ ;
  assign \new_Sorter100|0363_  = \new_Sorter100|0263_  & \new_Sorter100|0264_ ;
  assign \new_Sorter100|0364_  = \new_Sorter100|0263_  | \new_Sorter100|0264_ ;
  assign \new_Sorter100|0365_  = \new_Sorter100|0265_  & \new_Sorter100|0266_ ;
  assign \new_Sorter100|0366_  = \new_Sorter100|0265_  | \new_Sorter100|0266_ ;
  assign \new_Sorter100|0367_  = \new_Sorter100|0267_  & \new_Sorter100|0268_ ;
  assign \new_Sorter100|0368_  = \new_Sorter100|0267_  | \new_Sorter100|0268_ ;
  assign \new_Sorter100|0369_  = \new_Sorter100|0269_  & \new_Sorter100|0270_ ;
  assign \new_Sorter100|0370_  = \new_Sorter100|0269_  | \new_Sorter100|0270_ ;
  assign \new_Sorter100|0371_  = \new_Sorter100|0271_  & \new_Sorter100|0272_ ;
  assign \new_Sorter100|0372_  = \new_Sorter100|0271_  | \new_Sorter100|0272_ ;
  assign \new_Sorter100|0373_  = \new_Sorter100|0273_  & \new_Sorter100|0274_ ;
  assign \new_Sorter100|0374_  = \new_Sorter100|0273_  | \new_Sorter100|0274_ ;
  assign \new_Sorter100|0375_  = \new_Sorter100|0275_  & \new_Sorter100|0276_ ;
  assign \new_Sorter100|0376_  = \new_Sorter100|0275_  | \new_Sorter100|0276_ ;
  assign \new_Sorter100|0377_  = \new_Sorter100|0277_  & \new_Sorter100|0278_ ;
  assign \new_Sorter100|0378_  = \new_Sorter100|0277_  | \new_Sorter100|0278_ ;
  assign \new_Sorter100|0379_  = \new_Sorter100|0279_  & \new_Sorter100|0280_ ;
  assign \new_Sorter100|0380_  = \new_Sorter100|0279_  | \new_Sorter100|0280_ ;
  assign \new_Sorter100|0381_  = \new_Sorter100|0281_  & \new_Sorter100|0282_ ;
  assign \new_Sorter100|0382_  = \new_Sorter100|0281_  | \new_Sorter100|0282_ ;
  assign \new_Sorter100|0383_  = \new_Sorter100|0283_  & \new_Sorter100|0284_ ;
  assign \new_Sorter100|0384_  = \new_Sorter100|0283_  | \new_Sorter100|0284_ ;
  assign \new_Sorter100|0385_  = \new_Sorter100|0285_  & \new_Sorter100|0286_ ;
  assign \new_Sorter100|0386_  = \new_Sorter100|0285_  | \new_Sorter100|0286_ ;
  assign \new_Sorter100|0387_  = \new_Sorter100|0287_  & \new_Sorter100|0288_ ;
  assign \new_Sorter100|0388_  = \new_Sorter100|0287_  | \new_Sorter100|0288_ ;
  assign \new_Sorter100|0389_  = \new_Sorter100|0289_  & \new_Sorter100|0290_ ;
  assign \new_Sorter100|0390_  = \new_Sorter100|0289_  | \new_Sorter100|0290_ ;
  assign \new_Sorter100|0391_  = \new_Sorter100|0291_  & \new_Sorter100|0292_ ;
  assign \new_Sorter100|0392_  = \new_Sorter100|0291_  | \new_Sorter100|0292_ ;
  assign \new_Sorter100|0393_  = \new_Sorter100|0293_  & \new_Sorter100|0294_ ;
  assign \new_Sorter100|0394_  = \new_Sorter100|0293_  | \new_Sorter100|0294_ ;
  assign \new_Sorter100|0395_  = \new_Sorter100|0295_  & \new_Sorter100|0296_ ;
  assign \new_Sorter100|0396_  = \new_Sorter100|0295_  | \new_Sorter100|0296_ ;
  assign \new_Sorter100|0397_  = \new_Sorter100|0297_  & \new_Sorter100|0298_ ;
  assign \new_Sorter100|0398_  = \new_Sorter100|0297_  | \new_Sorter100|0298_ ;
  assign \new_Sorter100|0400_  = \new_Sorter100|0300_  & \new_Sorter100|0301_ ;
  assign \new_Sorter100|0401_  = \new_Sorter100|0300_  | \new_Sorter100|0301_ ;
  assign \new_Sorter100|0402_  = \new_Sorter100|0302_  & \new_Sorter100|0303_ ;
  assign \new_Sorter100|0403_  = \new_Sorter100|0302_  | \new_Sorter100|0303_ ;
  assign \new_Sorter100|0404_  = \new_Sorter100|0304_  & \new_Sorter100|0305_ ;
  assign \new_Sorter100|0405_  = \new_Sorter100|0304_  | \new_Sorter100|0305_ ;
  assign \new_Sorter100|0406_  = \new_Sorter100|0306_  & \new_Sorter100|0307_ ;
  assign \new_Sorter100|0407_  = \new_Sorter100|0306_  | \new_Sorter100|0307_ ;
  assign \new_Sorter100|0408_  = \new_Sorter100|0308_  & \new_Sorter100|0309_ ;
  assign \new_Sorter100|0409_  = \new_Sorter100|0308_  | \new_Sorter100|0309_ ;
  assign \new_Sorter100|0410_  = \new_Sorter100|0310_  & \new_Sorter100|0311_ ;
  assign \new_Sorter100|0411_  = \new_Sorter100|0310_  | \new_Sorter100|0311_ ;
  assign \new_Sorter100|0412_  = \new_Sorter100|0312_  & \new_Sorter100|0313_ ;
  assign \new_Sorter100|0413_  = \new_Sorter100|0312_  | \new_Sorter100|0313_ ;
  assign \new_Sorter100|0414_  = \new_Sorter100|0314_  & \new_Sorter100|0315_ ;
  assign \new_Sorter100|0415_  = \new_Sorter100|0314_  | \new_Sorter100|0315_ ;
  assign \new_Sorter100|0416_  = \new_Sorter100|0316_  & \new_Sorter100|0317_ ;
  assign \new_Sorter100|0417_  = \new_Sorter100|0316_  | \new_Sorter100|0317_ ;
  assign \new_Sorter100|0418_  = \new_Sorter100|0318_  & \new_Sorter100|0319_ ;
  assign \new_Sorter100|0419_  = \new_Sorter100|0318_  | \new_Sorter100|0319_ ;
  assign \new_Sorter100|0420_  = \new_Sorter100|0320_  & \new_Sorter100|0321_ ;
  assign \new_Sorter100|0421_  = \new_Sorter100|0320_  | \new_Sorter100|0321_ ;
  assign \new_Sorter100|0422_  = \new_Sorter100|0322_  & \new_Sorter100|0323_ ;
  assign \new_Sorter100|0423_  = \new_Sorter100|0322_  | \new_Sorter100|0323_ ;
  assign \new_Sorter100|0424_  = \new_Sorter100|0324_  & \new_Sorter100|0325_ ;
  assign \new_Sorter100|0425_  = \new_Sorter100|0324_  | \new_Sorter100|0325_ ;
  assign \new_Sorter100|0426_  = \new_Sorter100|0326_  & \new_Sorter100|0327_ ;
  assign \new_Sorter100|0427_  = \new_Sorter100|0326_  | \new_Sorter100|0327_ ;
  assign \new_Sorter100|0428_  = \new_Sorter100|0328_  & \new_Sorter100|0329_ ;
  assign \new_Sorter100|0429_  = \new_Sorter100|0328_  | \new_Sorter100|0329_ ;
  assign \new_Sorter100|0430_  = \new_Sorter100|0330_  & \new_Sorter100|0331_ ;
  assign \new_Sorter100|0431_  = \new_Sorter100|0330_  | \new_Sorter100|0331_ ;
  assign \new_Sorter100|0432_  = \new_Sorter100|0332_  & \new_Sorter100|0333_ ;
  assign \new_Sorter100|0433_  = \new_Sorter100|0332_  | \new_Sorter100|0333_ ;
  assign \new_Sorter100|0434_  = \new_Sorter100|0334_  & \new_Sorter100|0335_ ;
  assign \new_Sorter100|0435_  = \new_Sorter100|0334_  | \new_Sorter100|0335_ ;
  assign \new_Sorter100|0436_  = \new_Sorter100|0336_  & \new_Sorter100|0337_ ;
  assign \new_Sorter100|0437_  = \new_Sorter100|0336_  | \new_Sorter100|0337_ ;
  assign \new_Sorter100|0438_  = \new_Sorter100|0338_  & \new_Sorter100|0339_ ;
  assign \new_Sorter100|0439_  = \new_Sorter100|0338_  | \new_Sorter100|0339_ ;
  assign \new_Sorter100|0440_  = \new_Sorter100|0340_  & \new_Sorter100|0341_ ;
  assign \new_Sorter100|0441_  = \new_Sorter100|0340_  | \new_Sorter100|0341_ ;
  assign \new_Sorter100|0442_  = \new_Sorter100|0342_  & \new_Sorter100|0343_ ;
  assign \new_Sorter100|0443_  = \new_Sorter100|0342_  | \new_Sorter100|0343_ ;
  assign \new_Sorter100|0444_  = \new_Sorter100|0344_  & \new_Sorter100|0345_ ;
  assign \new_Sorter100|0445_  = \new_Sorter100|0344_  | \new_Sorter100|0345_ ;
  assign \new_Sorter100|0446_  = \new_Sorter100|0346_  & \new_Sorter100|0347_ ;
  assign \new_Sorter100|0447_  = \new_Sorter100|0346_  | \new_Sorter100|0347_ ;
  assign \new_Sorter100|0448_  = \new_Sorter100|0348_  & \new_Sorter100|0349_ ;
  assign \new_Sorter100|0449_  = \new_Sorter100|0348_  | \new_Sorter100|0349_ ;
  assign \new_Sorter100|0450_  = \new_Sorter100|0350_  & \new_Sorter100|0351_ ;
  assign \new_Sorter100|0451_  = \new_Sorter100|0350_  | \new_Sorter100|0351_ ;
  assign \new_Sorter100|0452_  = \new_Sorter100|0352_  & \new_Sorter100|0353_ ;
  assign \new_Sorter100|0453_  = \new_Sorter100|0352_  | \new_Sorter100|0353_ ;
  assign \new_Sorter100|0454_  = \new_Sorter100|0354_  & \new_Sorter100|0355_ ;
  assign \new_Sorter100|0455_  = \new_Sorter100|0354_  | \new_Sorter100|0355_ ;
  assign \new_Sorter100|0456_  = \new_Sorter100|0356_  & \new_Sorter100|0357_ ;
  assign \new_Sorter100|0457_  = \new_Sorter100|0356_  | \new_Sorter100|0357_ ;
  assign \new_Sorter100|0458_  = \new_Sorter100|0358_  & \new_Sorter100|0359_ ;
  assign \new_Sorter100|0459_  = \new_Sorter100|0358_  | \new_Sorter100|0359_ ;
  assign \new_Sorter100|0460_  = \new_Sorter100|0360_  & \new_Sorter100|0361_ ;
  assign \new_Sorter100|0461_  = \new_Sorter100|0360_  | \new_Sorter100|0361_ ;
  assign \new_Sorter100|0462_  = \new_Sorter100|0362_  & \new_Sorter100|0363_ ;
  assign \new_Sorter100|0463_  = \new_Sorter100|0362_  | \new_Sorter100|0363_ ;
  assign \new_Sorter100|0464_  = \new_Sorter100|0364_  & \new_Sorter100|0365_ ;
  assign \new_Sorter100|0465_  = \new_Sorter100|0364_  | \new_Sorter100|0365_ ;
  assign \new_Sorter100|0466_  = \new_Sorter100|0366_  & \new_Sorter100|0367_ ;
  assign \new_Sorter100|0467_  = \new_Sorter100|0366_  | \new_Sorter100|0367_ ;
  assign \new_Sorter100|0468_  = \new_Sorter100|0368_  & \new_Sorter100|0369_ ;
  assign \new_Sorter100|0469_  = \new_Sorter100|0368_  | \new_Sorter100|0369_ ;
  assign \new_Sorter100|0470_  = \new_Sorter100|0370_  & \new_Sorter100|0371_ ;
  assign \new_Sorter100|0471_  = \new_Sorter100|0370_  | \new_Sorter100|0371_ ;
  assign \new_Sorter100|0472_  = \new_Sorter100|0372_  & \new_Sorter100|0373_ ;
  assign \new_Sorter100|0473_  = \new_Sorter100|0372_  | \new_Sorter100|0373_ ;
  assign \new_Sorter100|0474_  = \new_Sorter100|0374_  & \new_Sorter100|0375_ ;
  assign \new_Sorter100|0475_  = \new_Sorter100|0374_  | \new_Sorter100|0375_ ;
  assign \new_Sorter100|0476_  = \new_Sorter100|0376_  & \new_Sorter100|0377_ ;
  assign \new_Sorter100|0477_  = \new_Sorter100|0376_  | \new_Sorter100|0377_ ;
  assign \new_Sorter100|0478_  = \new_Sorter100|0378_  & \new_Sorter100|0379_ ;
  assign \new_Sorter100|0479_  = \new_Sorter100|0378_  | \new_Sorter100|0379_ ;
  assign \new_Sorter100|0480_  = \new_Sorter100|0380_  & \new_Sorter100|0381_ ;
  assign \new_Sorter100|0481_  = \new_Sorter100|0380_  | \new_Sorter100|0381_ ;
  assign \new_Sorter100|0482_  = \new_Sorter100|0382_  & \new_Sorter100|0383_ ;
  assign \new_Sorter100|0483_  = \new_Sorter100|0382_  | \new_Sorter100|0383_ ;
  assign \new_Sorter100|0484_  = \new_Sorter100|0384_  & \new_Sorter100|0385_ ;
  assign \new_Sorter100|0485_  = \new_Sorter100|0384_  | \new_Sorter100|0385_ ;
  assign \new_Sorter100|0486_  = \new_Sorter100|0386_  & \new_Sorter100|0387_ ;
  assign \new_Sorter100|0487_  = \new_Sorter100|0386_  | \new_Sorter100|0387_ ;
  assign \new_Sorter100|0488_  = \new_Sorter100|0388_  & \new_Sorter100|0389_ ;
  assign \new_Sorter100|0489_  = \new_Sorter100|0388_  | \new_Sorter100|0389_ ;
  assign \new_Sorter100|0490_  = \new_Sorter100|0390_  & \new_Sorter100|0391_ ;
  assign \new_Sorter100|0491_  = \new_Sorter100|0390_  | \new_Sorter100|0391_ ;
  assign \new_Sorter100|0492_  = \new_Sorter100|0392_  & \new_Sorter100|0393_ ;
  assign \new_Sorter100|0493_  = \new_Sorter100|0392_  | \new_Sorter100|0393_ ;
  assign \new_Sorter100|0494_  = \new_Sorter100|0394_  & \new_Sorter100|0395_ ;
  assign \new_Sorter100|0495_  = \new_Sorter100|0394_  | \new_Sorter100|0395_ ;
  assign \new_Sorter100|0496_  = \new_Sorter100|0396_  & \new_Sorter100|0397_ ;
  assign \new_Sorter100|0497_  = \new_Sorter100|0396_  | \new_Sorter100|0397_ ;
  assign \new_Sorter100|0498_  = \new_Sorter100|0398_  & \new_Sorter100|0399_ ;
  assign \new_Sorter100|0499_  = \new_Sorter100|0398_  | \new_Sorter100|0399_ ;
  assign \new_Sorter100|0500_  = \new_Sorter100|0400_ ;
  assign \new_Sorter100|0599_  = \new_Sorter100|0499_ ;
  assign \new_Sorter100|0501_  = \new_Sorter100|0401_  & \new_Sorter100|0402_ ;
  assign \new_Sorter100|0502_  = \new_Sorter100|0401_  | \new_Sorter100|0402_ ;
  assign \new_Sorter100|0503_  = \new_Sorter100|0403_  & \new_Sorter100|0404_ ;
  assign \new_Sorter100|0504_  = \new_Sorter100|0403_  | \new_Sorter100|0404_ ;
  assign \new_Sorter100|0505_  = \new_Sorter100|0405_  & \new_Sorter100|0406_ ;
  assign \new_Sorter100|0506_  = \new_Sorter100|0405_  | \new_Sorter100|0406_ ;
  assign \new_Sorter100|0507_  = \new_Sorter100|0407_  & \new_Sorter100|0408_ ;
  assign \new_Sorter100|0508_  = \new_Sorter100|0407_  | \new_Sorter100|0408_ ;
  assign \new_Sorter100|0509_  = \new_Sorter100|0409_  & \new_Sorter100|0410_ ;
  assign \new_Sorter100|0510_  = \new_Sorter100|0409_  | \new_Sorter100|0410_ ;
  assign \new_Sorter100|0511_  = \new_Sorter100|0411_  & \new_Sorter100|0412_ ;
  assign \new_Sorter100|0512_  = \new_Sorter100|0411_  | \new_Sorter100|0412_ ;
  assign \new_Sorter100|0513_  = \new_Sorter100|0413_  & \new_Sorter100|0414_ ;
  assign \new_Sorter100|0514_  = \new_Sorter100|0413_  | \new_Sorter100|0414_ ;
  assign \new_Sorter100|0515_  = \new_Sorter100|0415_  & \new_Sorter100|0416_ ;
  assign \new_Sorter100|0516_  = \new_Sorter100|0415_  | \new_Sorter100|0416_ ;
  assign \new_Sorter100|0517_  = \new_Sorter100|0417_  & \new_Sorter100|0418_ ;
  assign \new_Sorter100|0518_  = \new_Sorter100|0417_  | \new_Sorter100|0418_ ;
  assign \new_Sorter100|0519_  = \new_Sorter100|0419_  & \new_Sorter100|0420_ ;
  assign \new_Sorter100|0520_  = \new_Sorter100|0419_  | \new_Sorter100|0420_ ;
  assign \new_Sorter100|0521_  = \new_Sorter100|0421_  & \new_Sorter100|0422_ ;
  assign \new_Sorter100|0522_  = \new_Sorter100|0421_  | \new_Sorter100|0422_ ;
  assign \new_Sorter100|0523_  = \new_Sorter100|0423_  & \new_Sorter100|0424_ ;
  assign \new_Sorter100|0524_  = \new_Sorter100|0423_  | \new_Sorter100|0424_ ;
  assign \new_Sorter100|0525_  = \new_Sorter100|0425_  & \new_Sorter100|0426_ ;
  assign \new_Sorter100|0526_  = \new_Sorter100|0425_  | \new_Sorter100|0426_ ;
  assign \new_Sorter100|0527_  = \new_Sorter100|0427_  & \new_Sorter100|0428_ ;
  assign \new_Sorter100|0528_  = \new_Sorter100|0427_  | \new_Sorter100|0428_ ;
  assign \new_Sorter100|0529_  = \new_Sorter100|0429_  & \new_Sorter100|0430_ ;
  assign \new_Sorter100|0530_  = \new_Sorter100|0429_  | \new_Sorter100|0430_ ;
  assign \new_Sorter100|0531_  = \new_Sorter100|0431_  & \new_Sorter100|0432_ ;
  assign \new_Sorter100|0532_  = \new_Sorter100|0431_  | \new_Sorter100|0432_ ;
  assign \new_Sorter100|0533_  = \new_Sorter100|0433_  & \new_Sorter100|0434_ ;
  assign \new_Sorter100|0534_  = \new_Sorter100|0433_  | \new_Sorter100|0434_ ;
  assign \new_Sorter100|0535_  = \new_Sorter100|0435_  & \new_Sorter100|0436_ ;
  assign \new_Sorter100|0536_  = \new_Sorter100|0435_  | \new_Sorter100|0436_ ;
  assign \new_Sorter100|0537_  = \new_Sorter100|0437_  & \new_Sorter100|0438_ ;
  assign \new_Sorter100|0538_  = \new_Sorter100|0437_  | \new_Sorter100|0438_ ;
  assign \new_Sorter100|0539_  = \new_Sorter100|0439_  & \new_Sorter100|0440_ ;
  assign \new_Sorter100|0540_  = \new_Sorter100|0439_  | \new_Sorter100|0440_ ;
  assign \new_Sorter100|0541_  = \new_Sorter100|0441_  & \new_Sorter100|0442_ ;
  assign \new_Sorter100|0542_  = \new_Sorter100|0441_  | \new_Sorter100|0442_ ;
  assign \new_Sorter100|0543_  = \new_Sorter100|0443_  & \new_Sorter100|0444_ ;
  assign \new_Sorter100|0544_  = \new_Sorter100|0443_  | \new_Sorter100|0444_ ;
  assign \new_Sorter100|0545_  = \new_Sorter100|0445_  & \new_Sorter100|0446_ ;
  assign \new_Sorter100|0546_  = \new_Sorter100|0445_  | \new_Sorter100|0446_ ;
  assign \new_Sorter100|0547_  = \new_Sorter100|0447_  & \new_Sorter100|0448_ ;
  assign \new_Sorter100|0548_  = \new_Sorter100|0447_  | \new_Sorter100|0448_ ;
  assign \new_Sorter100|0549_  = \new_Sorter100|0449_  & \new_Sorter100|0450_ ;
  assign \new_Sorter100|0550_  = \new_Sorter100|0449_  | \new_Sorter100|0450_ ;
  assign \new_Sorter100|0551_  = \new_Sorter100|0451_  & \new_Sorter100|0452_ ;
  assign \new_Sorter100|0552_  = \new_Sorter100|0451_  | \new_Sorter100|0452_ ;
  assign \new_Sorter100|0553_  = \new_Sorter100|0453_  & \new_Sorter100|0454_ ;
  assign \new_Sorter100|0554_  = \new_Sorter100|0453_  | \new_Sorter100|0454_ ;
  assign \new_Sorter100|0555_  = \new_Sorter100|0455_  & \new_Sorter100|0456_ ;
  assign \new_Sorter100|0556_  = \new_Sorter100|0455_  | \new_Sorter100|0456_ ;
  assign \new_Sorter100|0557_  = \new_Sorter100|0457_  & \new_Sorter100|0458_ ;
  assign \new_Sorter100|0558_  = \new_Sorter100|0457_  | \new_Sorter100|0458_ ;
  assign \new_Sorter100|0559_  = \new_Sorter100|0459_  & \new_Sorter100|0460_ ;
  assign \new_Sorter100|0560_  = \new_Sorter100|0459_  | \new_Sorter100|0460_ ;
  assign \new_Sorter100|0561_  = \new_Sorter100|0461_  & \new_Sorter100|0462_ ;
  assign \new_Sorter100|0562_  = \new_Sorter100|0461_  | \new_Sorter100|0462_ ;
  assign \new_Sorter100|0563_  = \new_Sorter100|0463_  & \new_Sorter100|0464_ ;
  assign \new_Sorter100|0564_  = \new_Sorter100|0463_  | \new_Sorter100|0464_ ;
  assign \new_Sorter100|0565_  = \new_Sorter100|0465_  & \new_Sorter100|0466_ ;
  assign \new_Sorter100|0566_  = \new_Sorter100|0465_  | \new_Sorter100|0466_ ;
  assign \new_Sorter100|0567_  = \new_Sorter100|0467_  & \new_Sorter100|0468_ ;
  assign \new_Sorter100|0568_  = \new_Sorter100|0467_  | \new_Sorter100|0468_ ;
  assign \new_Sorter100|0569_  = \new_Sorter100|0469_  & \new_Sorter100|0470_ ;
  assign \new_Sorter100|0570_  = \new_Sorter100|0469_  | \new_Sorter100|0470_ ;
  assign \new_Sorter100|0571_  = \new_Sorter100|0471_  & \new_Sorter100|0472_ ;
  assign \new_Sorter100|0572_  = \new_Sorter100|0471_  | \new_Sorter100|0472_ ;
  assign \new_Sorter100|0573_  = \new_Sorter100|0473_  & \new_Sorter100|0474_ ;
  assign \new_Sorter100|0574_  = \new_Sorter100|0473_  | \new_Sorter100|0474_ ;
  assign \new_Sorter100|0575_  = \new_Sorter100|0475_  & \new_Sorter100|0476_ ;
  assign \new_Sorter100|0576_  = \new_Sorter100|0475_  | \new_Sorter100|0476_ ;
  assign \new_Sorter100|0577_  = \new_Sorter100|0477_  & \new_Sorter100|0478_ ;
  assign \new_Sorter100|0578_  = \new_Sorter100|0477_  | \new_Sorter100|0478_ ;
  assign \new_Sorter100|0579_  = \new_Sorter100|0479_  & \new_Sorter100|0480_ ;
  assign \new_Sorter100|0580_  = \new_Sorter100|0479_  | \new_Sorter100|0480_ ;
  assign \new_Sorter100|0581_  = \new_Sorter100|0481_  & \new_Sorter100|0482_ ;
  assign \new_Sorter100|0582_  = \new_Sorter100|0481_  | \new_Sorter100|0482_ ;
  assign \new_Sorter100|0583_  = \new_Sorter100|0483_  & \new_Sorter100|0484_ ;
  assign \new_Sorter100|0584_  = \new_Sorter100|0483_  | \new_Sorter100|0484_ ;
  assign \new_Sorter100|0585_  = \new_Sorter100|0485_  & \new_Sorter100|0486_ ;
  assign \new_Sorter100|0586_  = \new_Sorter100|0485_  | \new_Sorter100|0486_ ;
  assign \new_Sorter100|0587_  = \new_Sorter100|0487_  & \new_Sorter100|0488_ ;
  assign \new_Sorter100|0588_  = \new_Sorter100|0487_  | \new_Sorter100|0488_ ;
  assign \new_Sorter100|0589_  = \new_Sorter100|0489_  & \new_Sorter100|0490_ ;
  assign \new_Sorter100|0590_  = \new_Sorter100|0489_  | \new_Sorter100|0490_ ;
  assign \new_Sorter100|0591_  = \new_Sorter100|0491_  & \new_Sorter100|0492_ ;
  assign \new_Sorter100|0592_  = \new_Sorter100|0491_  | \new_Sorter100|0492_ ;
  assign \new_Sorter100|0593_  = \new_Sorter100|0493_  & \new_Sorter100|0494_ ;
  assign \new_Sorter100|0594_  = \new_Sorter100|0493_  | \new_Sorter100|0494_ ;
  assign \new_Sorter100|0595_  = \new_Sorter100|0495_  & \new_Sorter100|0496_ ;
  assign \new_Sorter100|0596_  = \new_Sorter100|0495_  | \new_Sorter100|0496_ ;
  assign \new_Sorter100|0597_  = \new_Sorter100|0497_  & \new_Sorter100|0498_ ;
  assign \new_Sorter100|0598_  = \new_Sorter100|0497_  | \new_Sorter100|0498_ ;
  assign \new_Sorter100|0600_  = \new_Sorter100|0500_  & \new_Sorter100|0501_ ;
  assign \new_Sorter100|0601_  = \new_Sorter100|0500_  | \new_Sorter100|0501_ ;
  assign \new_Sorter100|0602_  = \new_Sorter100|0502_  & \new_Sorter100|0503_ ;
  assign \new_Sorter100|0603_  = \new_Sorter100|0502_  | \new_Sorter100|0503_ ;
  assign \new_Sorter100|0604_  = \new_Sorter100|0504_  & \new_Sorter100|0505_ ;
  assign \new_Sorter100|0605_  = \new_Sorter100|0504_  | \new_Sorter100|0505_ ;
  assign \new_Sorter100|0606_  = \new_Sorter100|0506_  & \new_Sorter100|0507_ ;
  assign \new_Sorter100|0607_  = \new_Sorter100|0506_  | \new_Sorter100|0507_ ;
  assign \new_Sorter100|0608_  = \new_Sorter100|0508_  & \new_Sorter100|0509_ ;
  assign \new_Sorter100|0609_  = \new_Sorter100|0508_  | \new_Sorter100|0509_ ;
  assign \new_Sorter100|0610_  = \new_Sorter100|0510_  & \new_Sorter100|0511_ ;
  assign \new_Sorter100|0611_  = \new_Sorter100|0510_  | \new_Sorter100|0511_ ;
  assign \new_Sorter100|0612_  = \new_Sorter100|0512_  & \new_Sorter100|0513_ ;
  assign \new_Sorter100|0613_  = \new_Sorter100|0512_  | \new_Sorter100|0513_ ;
  assign \new_Sorter100|0614_  = \new_Sorter100|0514_  & \new_Sorter100|0515_ ;
  assign \new_Sorter100|0615_  = \new_Sorter100|0514_  | \new_Sorter100|0515_ ;
  assign \new_Sorter100|0616_  = \new_Sorter100|0516_  & \new_Sorter100|0517_ ;
  assign \new_Sorter100|0617_  = \new_Sorter100|0516_  | \new_Sorter100|0517_ ;
  assign \new_Sorter100|0618_  = \new_Sorter100|0518_  & \new_Sorter100|0519_ ;
  assign \new_Sorter100|0619_  = \new_Sorter100|0518_  | \new_Sorter100|0519_ ;
  assign \new_Sorter100|0620_  = \new_Sorter100|0520_  & \new_Sorter100|0521_ ;
  assign \new_Sorter100|0621_  = \new_Sorter100|0520_  | \new_Sorter100|0521_ ;
  assign \new_Sorter100|0622_  = \new_Sorter100|0522_  & \new_Sorter100|0523_ ;
  assign \new_Sorter100|0623_  = \new_Sorter100|0522_  | \new_Sorter100|0523_ ;
  assign \new_Sorter100|0624_  = \new_Sorter100|0524_  & \new_Sorter100|0525_ ;
  assign \new_Sorter100|0625_  = \new_Sorter100|0524_  | \new_Sorter100|0525_ ;
  assign \new_Sorter100|0626_  = \new_Sorter100|0526_  & \new_Sorter100|0527_ ;
  assign \new_Sorter100|0627_  = \new_Sorter100|0526_  | \new_Sorter100|0527_ ;
  assign \new_Sorter100|0628_  = \new_Sorter100|0528_  & \new_Sorter100|0529_ ;
  assign \new_Sorter100|0629_  = \new_Sorter100|0528_  | \new_Sorter100|0529_ ;
  assign \new_Sorter100|0630_  = \new_Sorter100|0530_  & \new_Sorter100|0531_ ;
  assign \new_Sorter100|0631_  = \new_Sorter100|0530_  | \new_Sorter100|0531_ ;
  assign \new_Sorter100|0632_  = \new_Sorter100|0532_  & \new_Sorter100|0533_ ;
  assign \new_Sorter100|0633_  = \new_Sorter100|0532_  | \new_Sorter100|0533_ ;
  assign \new_Sorter100|0634_  = \new_Sorter100|0534_  & \new_Sorter100|0535_ ;
  assign \new_Sorter100|0635_  = \new_Sorter100|0534_  | \new_Sorter100|0535_ ;
  assign \new_Sorter100|0636_  = \new_Sorter100|0536_  & \new_Sorter100|0537_ ;
  assign \new_Sorter100|0637_  = \new_Sorter100|0536_  | \new_Sorter100|0537_ ;
  assign \new_Sorter100|0638_  = \new_Sorter100|0538_  & \new_Sorter100|0539_ ;
  assign \new_Sorter100|0639_  = \new_Sorter100|0538_  | \new_Sorter100|0539_ ;
  assign \new_Sorter100|0640_  = \new_Sorter100|0540_  & \new_Sorter100|0541_ ;
  assign \new_Sorter100|0641_  = \new_Sorter100|0540_  | \new_Sorter100|0541_ ;
  assign \new_Sorter100|0642_  = \new_Sorter100|0542_  & \new_Sorter100|0543_ ;
  assign \new_Sorter100|0643_  = \new_Sorter100|0542_  | \new_Sorter100|0543_ ;
  assign \new_Sorter100|0644_  = \new_Sorter100|0544_  & \new_Sorter100|0545_ ;
  assign \new_Sorter100|0645_  = \new_Sorter100|0544_  | \new_Sorter100|0545_ ;
  assign \new_Sorter100|0646_  = \new_Sorter100|0546_  & \new_Sorter100|0547_ ;
  assign \new_Sorter100|0647_  = \new_Sorter100|0546_  | \new_Sorter100|0547_ ;
  assign \new_Sorter100|0648_  = \new_Sorter100|0548_  & \new_Sorter100|0549_ ;
  assign \new_Sorter100|0649_  = \new_Sorter100|0548_  | \new_Sorter100|0549_ ;
  assign \new_Sorter100|0650_  = \new_Sorter100|0550_  & \new_Sorter100|0551_ ;
  assign \new_Sorter100|0651_  = \new_Sorter100|0550_  | \new_Sorter100|0551_ ;
  assign \new_Sorter100|0652_  = \new_Sorter100|0552_  & \new_Sorter100|0553_ ;
  assign \new_Sorter100|0653_  = \new_Sorter100|0552_  | \new_Sorter100|0553_ ;
  assign \new_Sorter100|0654_  = \new_Sorter100|0554_  & \new_Sorter100|0555_ ;
  assign \new_Sorter100|0655_  = \new_Sorter100|0554_  | \new_Sorter100|0555_ ;
  assign \new_Sorter100|0656_  = \new_Sorter100|0556_  & \new_Sorter100|0557_ ;
  assign \new_Sorter100|0657_  = \new_Sorter100|0556_  | \new_Sorter100|0557_ ;
  assign \new_Sorter100|0658_  = \new_Sorter100|0558_  & \new_Sorter100|0559_ ;
  assign \new_Sorter100|0659_  = \new_Sorter100|0558_  | \new_Sorter100|0559_ ;
  assign \new_Sorter100|0660_  = \new_Sorter100|0560_  & \new_Sorter100|0561_ ;
  assign \new_Sorter100|0661_  = \new_Sorter100|0560_  | \new_Sorter100|0561_ ;
  assign \new_Sorter100|0662_  = \new_Sorter100|0562_  & \new_Sorter100|0563_ ;
  assign \new_Sorter100|0663_  = \new_Sorter100|0562_  | \new_Sorter100|0563_ ;
  assign \new_Sorter100|0664_  = \new_Sorter100|0564_  & \new_Sorter100|0565_ ;
  assign \new_Sorter100|0665_  = \new_Sorter100|0564_  | \new_Sorter100|0565_ ;
  assign \new_Sorter100|0666_  = \new_Sorter100|0566_  & \new_Sorter100|0567_ ;
  assign \new_Sorter100|0667_  = \new_Sorter100|0566_  | \new_Sorter100|0567_ ;
  assign \new_Sorter100|0668_  = \new_Sorter100|0568_  & \new_Sorter100|0569_ ;
  assign \new_Sorter100|0669_  = \new_Sorter100|0568_  | \new_Sorter100|0569_ ;
  assign \new_Sorter100|0670_  = \new_Sorter100|0570_  & \new_Sorter100|0571_ ;
  assign \new_Sorter100|0671_  = \new_Sorter100|0570_  | \new_Sorter100|0571_ ;
  assign \new_Sorter100|0672_  = \new_Sorter100|0572_  & \new_Sorter100|0573_ ;
  assign \new_Sorter100|0673_  = \new_Sorter100|0572_  | \new_Sorter100|0573_ ;
  assign \new_Sorter100|0674_  = \new_Sorter100|0574_  & \new_Sorter100|0575_ ;
  assign \new_Sorter100|0675_  = \new_Sorter100|0574_  | \new_Sorter100|0575_ ;
  assign \new_Sorter100|0676_  = \new_Sorter100|0576_  & \new_Sorter100|0577_ ;
  assign \new_Sorter100|0677_  = \new_Sorter100|0576_  | \new_Sorter100|0577_ ;
  assign \new_Sorter100|0678_  = \new_Sorter100|0578_  & \new_Sorter100|0579_ ;
  assign \new_Sorter100|0679_  = \new_Sorter100|0578_  | \new_Sorter100|0579_ ;
  assign \new_Sorter100|0680_  = \new_Sorter100|0580_  & \new_Sorter100|0581_ ;
  assign \new_Sorter100|0681_  = \new_Sorter100|0580_  | \new_Sorter100|0581_ ;
  assign \new_Sorter100|0682_  = \new_Sorter100|0582_  & \new_Sorter100|0583_ ;
  assign \new_Sorter100|0683_  = \new_Sorter100|0582_  | \new_Sorter100|0583_ ;
  assign \new_Sorter100|0684_  = \new_Sorter100|0584_  & \new_Sorter100|0585_ ;
  assign \new_Sorter100|0685_  = \new_Sorter100|0584_  | \new_Sorter100|0585_ ;
  assign \new_Sorter100|0686_  = \new_Sorter100|0586_  & \new_Sorter100|0587_ ;
  assign \new_Sorter100|0687_  = \new_Sorter100|0586_  | \new_Sorter100|0587_ ;
  assign \new_Sorter100|0688_  = \new_Sorter100|0588_  & \new_Sorter100|0589_ ;
  assign \new_Sorter100|0689_  = \new_Sorter100|0588_  | \new_Sorter100|0589_ ;
  assign \new_Sorter100|0690_  = \new_Sorter100|0590_  & \new_Sorter100|0591_ ;
  assign \new_Sorter100|0691_  = \new_Sorter100|0590_  | \new_Sorter100|0591_ ;
  assign \new_Sorter100|0692_  = \new_Sorter100|0592_  & \new_Sorter100|0593_ ;
  assign \new_Sorter100|0693_  = \new_Sorter100|0592_  | \new_Sorter100|0593_ ;
  assign \new_Sorter100|0694_  = \new_Sorter100|0594_  & \new_Sorter100|0595_ ;
  assign \new_Sorter100|0695_  = \new_Sorter100|0594_  | \new_Sorter100|0595_ ;
  assign \new_Sorter100|0696_  = \new_Sorter100|0596_  & \new_Sorter100|0597_ ;
  assign \new_Sorter100|0697_  = \new_Sorter100|0596_  | \new_Sorter100|0597_ ;
  assign \new_Sorter100|0698_  = \new_Sorter100|0598_  & \new_Sorter100|0599_ ;
  assign \new_Sorter100|0699_  = \new_Sorter100|0598_  | \new_Sorter100|0599_ ;
  assign \new_Sorter100|0700_  = \new_Sorter100|0600_ ;
  assign \new_Sorter100|0799_  = \new_Sorter100|0699_ ;
  assign \new_Sorter100|0701_  = \new_Sorter100|0601_  & \new_Sorter100|0602_ ;
  assign \new_Sorter100|0702_  = \new_Sorter100|0601_  | \new_Sorter100|0602_ ;
  assign \new_Sorter100|0703_  = \new_Sorter100|0603_  & \new_Sorter100|0604_ ;
  assign \new_Sorter100|0704_  = \new_Sorter100|0603_  | \new_Sorter100|0604_ ;
  assign \new_Sorter100|0705_  = \new_Sorter100|0605_  & \new_Sorter100|0606_ ;
  assign \new_Sorter100|0706_  = \new_Sorter100|0605_  | \new_Sorter100|0606_ ;
  assign \new_Sorter100|0707_  = \new_Sorter100|0607_  & \new_Sorter100|0608_ ;
  assign \new_Sorter100|0708_  = \new_Sorter100|0607_  | \new_Sorter100|0608_ ;
  assign \new_Sorter100|0709_  = \new_Sorter100|0609_  & \new_Sorter100|0610_ ;
  assign \new_Sorter100|0710_  = \new_Sorter100|0609_  | \new_Sorter100|0610_ ;
  assign \new_Sorter100|0711_  = \new_Sorter100|0611_  & \new_Sorter100|0612_ ;
  assign \new_Sorter100|0712_  = \new_Sorter100|0611_  | \new_Sorter100|0612_ ;
  assign \new_Sorter100|0713_  = \new_Sorter100|0613_  & \new_Sorter100|0614_ ;
  assign \new_Sorter100|0714_  = \new_Sorter100|0613_  | \new_Sorter100|0614_ ;
  assign \new_Sorter100|0715_  = \new_Sorter100|0615_  & \new_Sorter100|0616_ ;
  assign \new_Sorter100|0716_  = \new_Sorter100|0615_  | \new_Sorter100|0616_ ;
  assign \new_Sorter100|0717_  = \new_Sorter100|0617_  & \new_Sorter100|0618_ ;
  assign \new_Sorter100|0718_  = \new_Sorter100|0617_  | \new_Sorter100|0618_ ;
  assign \new_Sorter100|0719_  = \new_Sorter100|0619_  & \new_Sorter100|0620_ ;
  assign \new_Sorter100|0720_  = \new_Sorter100|0619_  | \new_Sorter100|0620_ ;
  assign \new_Sorter100|0721_  = \new_Sorter100|0621_  & \new_Sorter100|0622_ ;
  assign \new_Sorter100|0722_  = \new_Sorter100|0621_  | \new_Sorter100|0622_ ;
  assign \new_Sorter100|0723_  = \new_Sorter100|0623_  & \new_Sorter100|0624_ ;
  assign \new_Sorter100|0724_  = \new_Sorter100|0623_  | \new_Sorter100|0624_ ;
  assign \new_Sorter100|0725_  = \new_Sorter100|0625_  & \new_Sorter100|0626_ ;
  assign \new_Sorter100|0726_  = \new_Sorter100|0625_  | \new_Sorter100|0626_ ;
  assign \new_Sorter100|0727_  = \new_Sorter100|0627_  & \new_Sorter100|0628_ ;
  assign \new_Sorter100|0728_  = \new_Sorter100|0627_  | \new_Sorter100|0628_ ;
  assign \new_Sorter100|0729_  = \new_Sorter100|0629_  & \new_Sorter100|0630_ ;
  assign \new_Sorter100|0730_  = \new_Sorter100|0629_  | \new_Sorter100|0630_ ;
  assign \new_Sorter100|0731_  = \new_Sorter100|0631_  & \new_Sorter100|0632_ ;
  assign \new_Sorter100|0732_  = \new_Sorter100|0631_  | \new_Sorter100|0632_ ;
  assign \new_Sorter100|0733_  = \new_Sorter100|0633_  & \new_Sorter100|0634_ ;
  assign \new_Sorter100|0734_  = \new_Sorter100|0633_  | \new_Sorter100|0634_ ;
  assign \new_Sorter100|0735_  = \new_Sorter100|0635_  & \new_Sorter100|0636_ ;
  assign \new_Sorter100|0736_  = \new_Sorter100|0635_  | \new_Sorter100|0636_ ;
  assign \new_Sorter100|0737_  = \new_Sorter100|0637_  & \new_Sorter100|0638_ ;
  assign \new_Sorter100|0738_  = \new_Sorter100|0637_  | \new_Sorter100|0638_ ;
  assign \new_Sorter100|0739_  = \new_Sorter100|0639_  & \new_Sorter100|0640_ ;
  assign \new_Sorter100|0740_  = \new_Sorter100|0639_  | \new_Sorter100|0640_ ;
  assign \new_Sorter100|0741_  = \new_Sorter100|0641_  & \new_Sorter100|0642_ ;
  assign \new_Sorter100|0742_  = \new_Sorter100|0641_  | \new_Sorter100|0642_ ;
  assign \new_Sorter100|0743_  = \new_Sorter100|0643_  & \new_Sorter100|0644_ ;
  assign \new_Sorter100|0744_  = \new_Sorter100|0643_  | \new_Sorter100|0644_ ;
  assign \new_Sorter100|0745_  = \new_Sorter100|0645_  & \new_Sorter100|0646_ ;
  assign \new_Sorter100|0746_  = \new_Sorter100|0645_  | \new_Sorter100|0646_ ;
  assign \new_Sorter100|0747_  = \new_Sorter100|0647_  & \new_Sorter100|0648_ ;
  assign \new_Sorter100|0748_  = \new_Sorter100|0647_  | \new_Sorter100|0648_ ;
  assign \new_Sorter100|0749_  = \new_Sorter100|0649_  & \new_Sorter100|0650_ ;
  assign \new_Sorter100|0750_  = \new_Sorter100|0649_  | \new_Sorter100|0650_ ;
  assign \new_Sorter100|0751_  = \new_Sorter100|0651_  & \new_Sorter100|0652_ ;
  assign \new_Sorter100|0752_  = \new_Sorter100|0651_  | \new_Sorter100|0652_ ;
  assign \new_Sorter100|0753_  = \new_Sorter100|0653_  & \new_Sorter100|0654_ ;
  assign \new_Sorter100|0754_  = \new_Sorter100|0653_  | \new_Sorter100|0654_ ;
  assign \new_Sorter100|0755_  = \new_Sorter100|0655_  & \new_Sorter100|0656_ ;
  assign \new_Sorter100|0756_  = \new_Sorter100|0655_  | \new_Sorter100|0656_ ;
  assign \new_Sorter100|0757_  = \new_Sorter100|0657_  & \new_Sorter100|0658_ ;
  assign \new_Sorter100|0758_  = \new_Sorter100|0657_  | \new_Sorter100|0658_ ;
  assign \new_Sorter100|0759_  = \new_Sorter100|0659_  & \new_Sorter100|0660_ ;
  assign \new_Sorter100|0760_  = \new_Sorter100|0659_  | \new_Sorter100|0660_ ;
  assign \new_Sorter100|0761_  = \new_Sorter100|0661_  & \new_Sorter100|0662_ ;
  assign \new_Sorter100|0762_  = \new_Sorter100|0661_  | \new_Sorter100|0662_ ;
  assign \new_Sorter100|0763_  = \new_Sorter100|0663_  & \new_Sorter100|0664_ ;
  assign \new_Sorter100|0764_  = \new_Sorter100|0663_  | \new_Sorter100|0664_ ;
  assign \new_Sorter100|0765_  = \new_Sorter100|0665_  & \new_Sorter100|0666_ ;
  assign \new_Sorter100|0766_  = \new_Sorter100|0665_  | \new_Sorter100|0666_ ;
  assign \new_Sorter100|0767_  = \new_Sorter100|0667_  & \new_Sorter100|0668_ ;
  assign \new_Sorter100|0768_  = \new_Sorter100|0667_  | \new_Sorter100|0668_ ;
  assign \new_Sorter100|0769_  = \new_Sorter100|0669_  & \new_Sorter100|0670_ ;
  assign \new_Sorter100|0770_  = \new_Sorter100|0669_  | \new_Sorter100|0670_ ;
  assign \new_Sorter100|0771_  = \new_Sorter100|0671_  & \new_Sorter100|0672_ ;
  assign \new_Sorter100|0772_  = \new_Sorter100|0671_  | \new_Sorter100|0672_ ;
  assign \new_Sorter100|0773_  = \new_Sorter100|0673_  & \new_Sorter100|0674_ ;
  assign \new_Sorter100|0774_  = \new_Sorter100|0673_  | \new_Sorter100|0674_ ;
  assign \new_Sorter100|0775_  = \new_Sorter100|0675_  & \new_Sorter100|0676_ ;
  assign \new_Sorter100|0776_  = \new_Sorter100|0675_  | \new_Sorter100|0676_ ;
  assign \new_Sorter100|0777_  = \new_Sorter100|0677_  & \new_Sorter100|0678_ ;
  assign \new_Sorter100|0778_  = \new_Sorter100|0677_  | \new_Sorter100|0678_ ;
  assign \new_Sorter100|0779_  = \new_Sorter100|0679_  & \new_Sorter100|0680_ ;
  assign \new_Sorter100|0780_  = \new_Sorter100|0679_  | \new_Sorter100|0680_ ;
  assign \new_Sorter100|0781_  = \new_Sorter100|0681_  & \new_Sorter100|0682_ ;
  assign \new_Sorter100|0782_  = \new_Sorter100|0681_  | \new_Sorter100|0682_ ;
  assign \new_Sorter100|0783_  = \new_Sorter100|0683_  & \new_Sorter100|0684_ ;
  assign \new_Sorter100|0784_  = \new_Sorter100|0683_  | \new_Sorter100|0684_ ;
  assign \new_Sorter100|0785_  = \new_Sorter100|0685_  & \new_Sorter100|0686_ ;
  assign \new_Sorter100|0786_  = \new_Sorter100|0685_  | \new_Sorter100|0686_ ;
  assign \new_Sorter100|0787_  = \new_Sorter100|0687_  & \new_Sorter100|0688_ ;
  assign \new_Sorter100|0788_  = \new_Sorter100|0687_  | \new_Sorter100|0688_ ;
  assign \new_Sorter100|0789_  = \new_Sorter100|0689_  & \new_Sorter100|0690_ ;
  assign \new_Sorter100|0790_  = \new_Sorter100|0689_  | \new_Sorter100|0690_ ;
  assign \new_Sorter100|0791_  = \new_Sorter100|0691_  & \new_Sorter100|0692_ ;
  assign \new_Sorter100|0792_  = \new_Sorter100|0691_  | \new_Sorter100|0692_ ;
  assign \new_Sorter100|0793_  = \new_Sorter100|0693_  & \new_Sorter100|0694_ ;
  assign \new_Sorter100|0794_  = \new_Sorter100|0693_  | \new_Sorter100|0694_ ;
  assign \new_Sorter100|0795_  = \new_Sorter100|0695_  & \new_Sorter100|0696_ ;
  assign \new_Sorter100|0796_  = \new_Sorter100|0695_  | \new_Sorter100|0696_ ;
  assign \new_Sorter100|0797_  = \new_Sorter100|0697_  & \new_Sorter100|0698_ ;
  assign \new_Sorter100|0798_  = \new_Sorter100|0697_  | \new_Sorter100|0698_ ;
  assign \new_Sorter100|0800_  = \new_Sorter100|0700_  & \new_Sorter100|0701_ ;
  assign \new_Sorter100|0801_  = \new_Sorter100|0700_  | \new_Sorter100|0701_ ;
  assign \new_Sorter100|0802_  = \new_Sorter100|0702_  & \new_Sorter100|0703_ ;
  assign \new_Sorter100|0803_  = \new_Sorter100|0702_  | \new_Sorter100|0703_ ;
  assign \new_Sorter100|0804_  = \new_Sorter100|0704_  & \new_Sorter100|0705_ ;
  assign \new_Sorter100|0805_  = \new_Sorter100|0704_  | \new_Sorter100|0705_ ;
  assign \new_Sorter100|0806_  = \new_Sorter100|0706_  & \new_Sorter100|0707_ ;
  assign \new_Sorter100|0807_  = \new_Sorter100|0706_  | \new_Sorter100|0707_ ;
  assign \new_Sorter100|0808_  = \new_Sorter100|0708_  & \new_Sorter100|0709_ ;
  assign \new_Sorter100|0809_  = \new_Sorter100|0708_  | \new_Sorter100|0709_ ;
  assign \new_Sorter100|0810_  = \new_Sorter100|0710_  & \new_Sorter100|0711_ ;
  assign \new_Sorter100|0811_  = \new_Sorter100|0710_  | \new_Sorter100|0711_ ;
  assign \new_Sorter100|0812_  = \new_Sorter100|0712_  & \new_Sorter100|0713_ ;
  assign \new_Sorter100|0813_  = \new_Sorter100|0712_  | \new_Sorter100|0713_ ;
  assign \new_Sorter100|0814_  = \new_Sorter100|0714_  & \new_Sorter100|0715_ ;
  assign \new_Sorter100|0815_  = \new_Sorter100|0714_  | \new_Sorter100|0715_ ;
  assign \new_Sorter100|0816_  = \new_Sorter100|0716_  & \new_Sorter100|0717_ ;
  assign \new_Sorter100|0817_  = \new_Sorter100|0716_  | \new_Sorter100|0717_ ;
  assign \new_Sorter100|0818_  = \new_Sorter100|0718_  & \new_Sorter100|0719_ ;
  assign \new_Sorter100|0819_  = \new_Sorter100|0718_  | \new_Sorter100|0719_ ;
  assign \new_Sorter100|0820_  = \new_Sorter100|0720_  & \new_Sorter100|0721_ ;
  assign \new_Sorter100|0821_  = \new_Sorter100|0720_  | \new_Sorter100|0721_ ;
  assign \new_Sorter100|0822_  = \new_Sorter100|0722_  & \new_Sorter100|0723_ ;
  assign \new_Sorter100|0823_  = \new_Sorter100|0722_  | \new_Sorter100|0723_ ;
  assign \new_Sorter100|0824_  = \new_Sorter100|0724_  & \new_Sorter100|0725_ ;
  assign \new_Sorter100|0825_  = \new_Sorter100|0724_  | \new_Sorter100|0725_ ;
  assign \new_Sorter100|0826_  = \new_Sorter100|0726_  & \new_Sorter100|0727_ ;
  assign \new_Sorter100|0827_  = \new_Sorter100|0726_  | \new_Sorter100|0727_ ;
  assign \new_Sorter100|0828_  = \new_Sorter100|0728_  & \new_Sorter100|0729_ ;
  assign \new_Sorter100|0829_  = \new_Sorter100|0728_  | \new_Sorter100|0729_ ;
  assign \new_Sorter100|0830_  = \new_Sorter100|0730_  & \new_Sorter100|0731_ ;
  assign \new_Sorter100|0831_  = \new_Sorter100|0730_  | \new_Sorter100|0731_ ;
  assign \new_Sorter100|0832_  = \new_Sorter100|0732_  & \new_Sorter100|0733_ ;
  assign \new_Sorter100|0833_  = \new_Sorter100|0732_  | \new_Sorter100|0733_ ;
  assign \new_Sorter100|0834_  = \new_Sorter100|0734_  & \new_Sorter100|0735_ ;
  assign \new_Sorter100|0835_  = \new_Sorter100|0734_  | \new_Sorter100|0735_ ;
  assign \new_Sorter100|0836_  = \new_Sorter100|0736_  & \new_Sorter100|0737_ ;
  assign \new_Sorter100|0837_  = \new_Sorter100|0736_  | \new_Sorter100|0737_ ;
  assign \new_Sorter100|0838_  = \new_Sorter100|0738_  & \new_Sorter100|0739_ ;
  assign \new_Sorter100|0839_  = \new_Sorter100|0738_  | \new_Sorter100|0739_ ;
  assign \new_Sorter100|0840_  = \new_Sorter100|0740_  & \new_Sorter100|0741_ ;
  assign \new_Sorter100|0841_  = \new_Sorter100|0740_  | \new_Sorter100|0741_ ;
  assign \new_Sorter100|0842_  = \new_Sorter100|0742_  & \new_Sorter100|0743_ ;
  assign \new_Sorter100|0843_  = \new_Sorter100|0742_  | \new_Sorter100|0743_ ;
  assign \new_Sorter100|0844_  = \new_Sorter100|0744_  & \new_Sorter100|0745_ ;
  assign \new_Sorter100|0845_  = \new_Sorter100|0744_  | \new_Sorter100|0745_ ;
  assign \new_Sorter100|0846_  = \new_Sorter100|0746_  & \new_Sorter100|0747_ ;
  assign \new_Sorter100|0847_  = \new_Sorter100|0746_  | \new_Sorter100|0747_ ;
  assign \new_Sorter100|0848_  = \new_Sorter100|0748_  & \new_Sorter100|0749_ ;
  assign \new_Sorter100|0849_  = \new_Sorter100|0748_  | \new_Sorter100|0749_ ;
  assign \new_Sorter100|0850_  = \new_Sorter100|0750_  & \new_Sorter100|0751_ ;
  assign \new_Sorter100|0851_  = \new_Sorter100|0750_  | \new_Sorter100|0751_ ;
  assign \new_Sorter100|0852_  = \new_Sorter100|0752_  & \new_Sorter100|0753_ ;
  assign \new_Sorter100|0853_  = \new_Sorter100|0752_  | \new_Sorter100|0753_ ;
  assign \new_Sorter100|0854_  = \new_Sorter100|0754_  & \new_Sorter100|0755_ ;
  assign \new_Sorter100|0855_  = \new_Sorter100|0754_  | \new_Sorter100|0755_ ;
  assign \new_Sorter100|0856_  = \new_Sorter100|0756_  & \new_Sorter100|0757_ ;
  assign \new_Sorter100|0857_  = \new_Sorter100|0756_  | \new_Sorter100|0757_ ;
  assign \new_Sorter100|0858_  = \new_Sorter100|0758_  & \new_Sorter100|0759_ ;
  assign \new_Sorter100|0859_  = \new_Sorter100|0758_  | \new_Sorter100|0759_ ;
  assign \new_Sorter100|0860_  = \new_Sorter100|0760_  & \new_Sorter100|0761_ ;
  assign \new_Sorter100|0861_  = \new_Sorter100|0760_  | \new_Sorter100|0761_ ;
  assign \new_Sorter100|0862_  = \new_Sorter100|0762_  & \new_Sorter100|0763_ ;
  assign \new_Sorter100|0863_  = \new_Sorter100|0762_  | \new_Sorter100|0763_ ;
  assign \new_Sorter100|0864_  = \new_Sorter100|0764_  & \new_Sorter100|0765_ ;
  assign \new_Sorter100|0865_  = \new_Sorter100|0764_  | \new_Sorter100|0765_ ;
  assign \new_Sorter100|0866_  = \new_Sorter100|0766_  & \new_Sorter100|0767_ ;
  assign \new_Sorter100|0867_  = \new_Sorter100|0766_  | \new_Sorter100|0767_ ;
  assign \new_Sorter100|0868_  = \new_Sorter100|0768_  & \new_Sorter100|0769_ ;
  assign \new_Sorter100|0869_  = \new_Sorter100|0768_  | \new_Sorter100|0769_ ;
  assign \new_Sorter100|0870_  = \new_Sorter100|0770_  & \new_Sorter100|0771_ ;
  assign \new_Sorter100|0871_  = \new_Sorter100|0770_  | \new_Sorter100|0771_ ;
  assign \new_Sorter100|0872_  = \new_Sorter100|0772_  & \new_Sorter100|0773_ ;
  assign \new_Sorter100|0873_  = \new_Sorter100|0772_  | \new_Sorter100|0773_ ;
  assign \new_Sorter100|0874_  = \new_Sorter100|0774_  & \new_Sorter100|0775_ ;
  assign \new_Sorter100|0875_  = \new_Sorter100|0774_  | \new_Sorter100|0775_ ;
  assign \new_Sorter100|0876_  = \new_Sorter100|0776_  & \new_Sorter100|0777_ ;
  assign \new_Sorter100|0877_  = \new_Sorter100|0776_  | \new_Sorter100|0777_ ;
  assign \new_Sorter100|0878_  = \new_Sorter100|0778_  & \new_Sorter100|0779_ ;
  assign \new_Sorter100|0879_  = \new_Sorter100|0778_  | \new_Sorter100|0779_ ;
  assign \new_Sorter100|0880_  = \new_Sorter100|0780_  & \new_Sorter100|0781_ ;
  assign \new_Sorter100|0881_  = \new_Sorter100|0780_  | \new_Sorter100|0781_ ;
  assign \new_Sorter100|0882_  = \new_Sorter100|0782_  & \new_Sorter100|0783_ ;
  assign \new_Sorter100|0883_  = \new_Sorter100|0782_  | \new_Sorter100|0783_ ;
  assign \new_Sorter100|0884_  = \new_Sorter100|0784_  & \new_Sorter100|0785_ ;
  assign \new_Sorter100|0885_  = \new_Sorter100|0784_  | \new_Sorter100|0785_ ;
  assign \new_Sorter100|0886_  = \new_Sorter100|0786_  & \new_Sorter100|0787_ ;
  assign \new_Sorter100|0887_  = \new_Sorter100|0786_  | \new_Sorter100|0787_ ;
  assign \new_Sorter100|0888_  = \new_Sorter100|0788_  & \new_Sorter100|0789_ ;
  assign \new_Sorter100|0889_  = \new_Sorter100|0788_  | \new_Sorter100|0789_ ;
  assign \new_Sorter100|0890_  = \new_Sorter100|0790_  & \new_Sorter100|0791_ ;
  assign \new_Sorter100|0891_  = \new_Sorter100|0790_  | \new_Sorter100|0791_ ;
  assign \new_Sorter100|0892_  = \new_Sorter100|0792_  & \new_Sorter100|0793_ ;
  assign \new_Sorter100|0893_  = \new_Sorter100|0792_  | \new_Sorter100|0793_ ;
  assign \new_Sorter100|0894_  = \new_Sorter100|0794_  & \new_Sorter100|0795_ ;
  assign \new_Sorter100|0895_  = \new_Sorter100|0794_  | \new_Sorter100|0795_ ;
  assign \new_Sorter100|0896_  = \new_Sorter100|0796_  & \new_Sorter100|0797_ ;
  assign \new_Sorter100|0897_  = \new_Sorter100|0796_  | \new_Sorter100|0797_ ;
  assign \new_Sorter100|0898_  = \new_Sorter100|0798_  & \new_Sorter100|0799_ ;
  assign \new_Sorter100|0899_  = \new_Sorter100|0798_  | \new_Sorter100|0799_ ;
  assign \new_Sorter100|0900_  = \new_Sorter100|0800_ ;
  assign \new_Sorter100|0999_  = \new_Sorter100|0899_ ;
  assign \new_Sorter100|0901_  = \new_Sorter100|0801_  & \new_Sorter100|0802_ ;
  assign \new_Sorter100|0902_  = \new_Sorter100|0801_  | \new_Sorter100|0802_ ;
  assign \new_Sorter100|0903_  = \new_Sorter100|0803_  & \new_Sorter100|0804_ ;
  assign \new_Sorter100|0904_  = \new_Sorter100|0803_  | \new_Sorter100|0804_ ;
  assign \new_Sorter100|0905_  = \new_Sorter100|0805_  & \new_Sorter100|0806_ ;
  assign \new_Sorter100|0906_  = \new_Sorter100|0805_  | \new_Sorter100|0806_ ;
  assign \new_Sorter100|0907_  = \new_Sorter100|0807_  & \new_Sorter100|0808_ ;
  assign \new_Sorter100|0908_  = \new_Sorter100|0807_  | \new_Sorter100|0808_ ;
  assign \new_Sorter100|0909_  = \new_Sorter100|0809_  & \new_Sorter100|0810_ ;
  assign \new_Sorter100|0910_  = \new_Sorter100|0809_  | \new_Sorter100|0810_ ;
  assign \new_Sorter100|0911_  = \new_Sorter100|0811_  & \new_Sorter100|0812_ ;
  assign \new_Sorter100|0912_  = \new_Sorter100|0811_  | \new_Sorter100|0812_ ;
  assign \new_Sorter100|0913_  = \new_Sorter100|0813_  & \new_Sorter100|0814_ ;
  assign \new_Sorter100|0914_  = \new_Sorter100|0813_  | \new_Sorter100|0814_ ;
  assign \new_Sorter100|0915_  = \new_Sorter100|0815_  & \new_Sorter100|0816_ ;
  assign \new_Sorter100|0916_  = \new_Sorter100|0815_  | \new_Sorter100|0816_ ;
  assign \new_Sorter100|0917_  = \new_Sorter100|0817_  & \new_Sorter100|0818_ ;
  assign \new_Sorter100|0918_  = \new_Sorter100|0817_  | \new_Sorter100|0818_ ;
  assign \new_Sorter100|0919_  = \new_Sorter100|0819_  & \new_Sorter100|0820_ ;
  assign \new_Sorter100|0920_  = \new_Sorter100|0819_  | \new_Sorter100|0820_ ;
  assign \new_Sorter100|0921_  = \new_Sorter100|0821_  & \new_Sorter100|0822_ ;
  assign \new_Sorter100|0922_  = \new_Sorter100|0821_  | \new_Sorter100|0822_ ;
  assign \new_Sorter100|0923_  = \new_Sorter100|0823_  & \new_Sorter100|0824_ ;
  assign \new_Sorter100|0924_  = \new_Sorter100|0823_  | \new_Sorter100|0824_ ;
  assign \new_Sorter100|0925_  = \new_Sorter100|0825_  & \new_Sorter100|0826_ ;
  assign \new_Sorter100|0926_  = \new_Sorter100|0825_  | \new_Sorter100|0826_ ;
  assign \new_Sorter100|0927_  = \new_Sorter100|0827_  & \new_Sorter100|0828_ ;
  assign \new_Sorter100|0928_  = \new_Sorter100|0827_  | \new_Sorter100|0828_ ;
  assign \new_Sorter100|0929_  = \new_Sorter100|0829_  & \new_Sorter100|0830_ ;
  assign \new_Sorter100|0930_  = \new_Sorter100|0829_  | \new_Sorter100|0830_ ;
  assign \new_Sorter100|0931_  = \new_Sorter100|0831_  & \new_Sorter100|0832_ ;
  assign \new_Sorter100|0932_  = \new_Sorter100|0831_  | \new_Sorter100|0832_ ;
  assign \new_Sorter100|0933_  = \new_Sorter100|0833_  & \new_Sorter100|0834_ ;
  assign \new_Sorter100|0934_  = \new_Sorter100|0833_  | \new_Sorter100|0834_ ;
  assign \new_Sorter100|0935_  = \new_Sorter100|0835_  & \new_Sorter100|0836_ ;
  assign \new_Sorter100|0936_  = \new_Sorter100|0835_  | \new_Sorter100|0836_ ;
  assign \new_Sorter100|0937_  = \new_Sorter100|0837_  & \new_Sorter100|0838_ ;
  assign \new_Sorter100|0938_  = \new_Sorter100|0837_  | \new_Sorter100|0838_ ;
  assign \new_Sorter100|0939_  = \new_Sorter100|0839_  & \new_Sorter100|0840_ ;
  assign \new_Sorter100|0940_  = \new_Sorter100|0839_  | \new_Sorter100|0840_ ;
  assign \new_Sorter100|0941_  = \new_Sorter100|0841_  & \new_Sorter100|0842_ ;
  assign \new_Sorter100|0942_  = \new_Sorter100|0841_  | \new_Sorter100|0842_ ;
  assign \new_Sorter100|0943_  = \new_Sorter100|0843_  & \new_Sorter100|0844_ ;
  assign \new_Sorter100|0944_  = \new_Sorter100|0843_  | \new_Sorter100|0844_ ;
  assign \new_Sorter100|0945_  = \new_Sorter100|0845_  & \new_Sorter100|0846_ ;
  assign \new_Sorter100|0946_  = \new_Sorter100|0845_  | \new_Sorter100|0846_ ;
  assign \new_Sorter100|0947_  = \new_Sorter100|0847_  & \new_Sorter100|0848_ ;
  assign \new_Sorter100|0948_  = \new_Sorter100|0847_  | \new_Sorter100|0848_ ;
  assign \new_Sorter100|0949_  = \new_Sorter100|0849_  & \new_Sorter100|0850_ ;
  assign \new_Sorter100|0950_  = \new_Sorter100|0849_  | \new_Sorter100|0850_ ;
  assign \new_Sorter100|0951_  = \new_Sorter100|0851_  & \new_Sorter100|0852_ ;
  assign \new_Sorter100|0952_  = \new_Sorter100|0851_  | \new_Sorter100|0852_ ;
  assign \new_Sorter100|0953_  = \new_Sorter100|0853_  & \new_Sorter100|0854_ ;
  assign \new_Sorter100|0954_  = \new_Sorter100|0853_  | \new_Sorter100|0854_ ;
  assign \new_Sorter100|0955_  = \new_Sorter100|0855_  & \new_Sorter100|0856_ ;
  assign \new_Sorter100|0956_  = \new_Sorter100|0855_  | \new_Sorter100|0856_ ;
  assign \new_Sorter100|0957_  = \new_Sorter100|0857_  & \new_Sorter100|0858_ ;
  assign \new_Sorter100|0958_  = \new_Sorter100|0857_  | \new_Sorter100|0858_ ;
  assign \new_Sorter100|0959_  = \new_Sorter100|0859_  & \new_Sorter100|0860_ ;
  assign \new_Sorter100|0960_  = \new_Sorter100|0859_  | \new_Sorter100|0860_ ;
  assign \new_Sorter100|0961_  = \new_Sorter100|0861_  & \new_Sorter100|0862_ ;
  assign \new_Sorter100|0962_  = \new_Sorter100|0861_  | \new_Sorter100|0862_ ;
  assign \new_Sorter100|0963_  = \new_Sorter100|0863_  & \new_Sorter100|0864_ ;
  assign \new_Sorter100|0964_  = \new_Sorter100|0863_  | \new_Sorter100|0864_ ;
  assign \new_Sorter100|0965_  = \new_Sorter100|0865_  & \new_Sorter100|0866_ ;
  assign \new_Sorter100|0966_  = \new_Sorter100|0865_  | \new_Sorter100|0866_ ;
  assign \new_Sorter100|0967_  = \new_Sorter100|0867_  & \new_Sorter100|0868_ ;
  assign \new_Sorter100|0968_  = \new_Sorter100|0867_  | \new_Sorter100|0868_ ;
  assign \new_Sorter100|0969_  = \new_Sorter100|0869_  & \new_Sorter100|0870_ ;
  assign \new_Sorter100|0970_  = \new_Sorter100|0869_  | \new_Sorter100|0870_ ;
  assign \new_Sorter100|0971_  = \new_Sorter100|0871_  & \new_Sorter100|0872_ ;
  assign \new_Sorter100|0972_  = \new_Sorter100|0871_  | \new_Sorter100|0872_ ;
  assign \new_Sorter100|0973_  = \new_Sorter100|0873_  & \new_Sorter100|0874_ ;
  assign \new_Sorter100|0974_  = \new_Sorter100|0873_  | \new_Sorter100|0874_ ;
  assign \new_Sorter100|0975_  = \new_Sorter100|0875_  & \new_Sorter100|0876_ ;
  assign \new_Sorter100|0976_  = \new_Sorter100|0875_  | \new_Sorter100|0876_ ;
  assign \new_Sorter100|0977_  = \new_Sorter100|0877_  & \new_Sorter100|0878_ ;
  assign \new_Sorter100|0978_  = \new_Sorter100|0877_  | \new_Sorter100|0878_ ;
  assign \new_Sorter100|0979_  = \new_Sorter100|0879_  & \new_Sorter100|0880_ ;
  assign \new_Sorter100|0980_  = \new_Sorter100|0879_  | \new_Sorter100|0880_ ;
  assign \new_Sorter100|0981_  = \new_Sorter100|0881_  & \new_Sorter100|0882_ ;
  assign \new_Sorter100|0982_  = \new_Sorter100|0881_  | \new_Sorter100|0882_ ;
  assign \new_Sorter100|0983_  = \new_Sorter100|0883_  & \new_Sorter100|0884_ ;
  assign \new_Sorter100|0984_  = \new_Sorter100|0883_  | \new_Sorter100|0884_ ;
  assign \new_Sorter100|0985_  = \new_Sorter100|0885_  & \new_Sorter100|0886_ ;
  assign \new_Sorter100|0986_  = \new_Sorter100|0885_  | \new_Sorter100|0886_ ;
  assign \new_Sorter100|0987_  = \new_Sorter100|0887_  & \new_Sorter100|0888_ ;
  assign \new_Sorter100|0988_  = \new_Sorter100|0887_  | \new_Sorter100|0888_ ;
  assign \new_Sorter100|0989_  = \new_Sorter100|0889_  & \new_Sorter100|0890_ ;
  assign \new_Sorter100|0990_  = \new_Sorter100|0889_  | \new_Sorter100|0890_ ;
  assign \new_Sorter100|0991_  = \new_Sorter100|0891_  & \new_Sorter100|0892_ ;
  assign \new_Sorter100|0992_  = \new_Sorter100|0891_  | \new_Sorter100|0892_ ;
  assign \new_Sorter100|0993_  = \new_Sorter100|0893_  & \new_Sorter100|0894_ ;
  assign \new_Sorter100|0994_  = \new_Sorter100|0893_  | \new_Sorter100|0894_ ;
  assign \new_Sorter100|0995_  = \new_Sorter100|0895_  & \new_Sorter100|0896_ ;
  assign \new_Sorter100|0996_  = \new_Sorter100|0895_  | \new_Sorter100|0896_ ;
  assign \new_Sorter100|0997_  = \new_Sorter100|0897_  & \new_Sorter100|0898_ ;
  assign \new_Sorter100|0998_  = \new_Sorter100|0897_  | \new_Sorter100|0898_ ;
  assign \new_Sorter100|1000_  = \new_Sorter100|0900_  & \new_Sorter100|0901_ ;
  assign \new_Sorter100|1001_  = \new_Sorter100|0900_  | \new_Sorter100|0901_ ;
  assign \new_Sorter100|1002_  = \new_Sorter100|0902_  & \new_Sorter100|0903_ ;
  assign \new_Sorter100|1003_  = \new_Sorter100|0902_  | \new_Sorter100|0903_ ;
  assign \new_Sorter100|1004_  = \new_Sorter100|0904_  & \new_Sorter100|0905_ ;
  assign \new_Sorter100|1005_  = \new_Sorter100|0904_  | \new_Sorter100|0905_ ;
  assign \new_Sorter100|1006_  = \new_Sorter100|0906_  & \new_Sorter100|0907_ ;
  assign \new_Sorter100|1007_  = \new_Sorter100|0906_  | \new_Sorter100|0907_ ;
  assign \new_Sorter100|1008_  = \new_Sorter100|0908_  & \new_Sorter100|0909_ ;
  assign \new_Sorter100|1009_  = \new_Sorter100|0908_  | \new_Sorter100|0909_ ;
  assign \new_Sorter100|1010_  = \new_Sorter100|0910_  & \new_Sorter100|0911_ ;
  assign \new_Sorter100|1011_  = \new_Sorter100|0910_  | \new_Sorter100|0911_ ;
  assign \new_Sorter100|1012_  = \new_Sorter100|0912_  & \new_Sorter100|0913_ ;
  assign \new_Sorter100|1013_  = \new_Sorter100|0912_  | \new_Sorter100|0913_ ;
  assign \new_Sorter100|1014_  = \new_Sorter100|0914_  & \new_Sorter100|0915_ ;
  assign \new_Sorter100|1015_  = \new_Sorter100|0914_  | \new_Sorter100|0915_ ;
  assign \new_Sorter100|1016_  = \new_Sorter100|0916_  & \new_Sorter100|0917_ ;
  assign \new_Sorter100|1017_  = \new_Sorter100|0916_  | \new_Sorter100|0917_ ;
  assign \new_Sorter100|1018_  = \new_Sorter100|0918_  & \new_Sorter100|0919_ ;
  assign \new_Sorter100|1019_  = \new_Sorter100|0918_  | \new_Sorter100|0919_ ;
  assign \new_Sorter100|1020_  = \new_Sorter100|0920_  & \new_Sorter100|0921_ ;
  assign \new_Sorter100|1021_  = \new_Sorter100|0920_  | \new_Sorter100|0921_ ;
  assign \new_Sorter100|1022_  = \new_Sorter100|0922_  & \new_Sorter100|0923_ ;
  assign \new_Sorter100|1023_  = \new_Sorter100|0922_  | \new_Sorter100|0923_ ;
  assign \new_Sorter100|1024_  = \new_Sorter100|0924_  & \new_Sorter100|0925_ ;
  assign \new_Sorter100|1025_  = \new_Sorter100|0924_  | \new_Sorter100|0925_ ;
  assign \new_Sorter100|1026_  = \new_Sorter100|0926_  & \new_Sorter100|0927_ ;
  assign \new_Sorter100|1027_  = \new_Sorter100|0926_  | \new_Sorter100|0927_ ;
  assign \new_Sorter100|1028_  = \new_Sorter100|0928_  & \new_Sorter100|0929_ ;
  assign \new_Sorter100|1029_  = \new_Sorter100|0928_  | \new_Sorter100|0929_ ;
  assign \new_Sorter100|1030_  = \new_Sorter100|0930_  & \new_Sorter100|0931_ ;
  assign \new_Sorter100|1031_  = \new_Sorter100|0930_  | \new_Sorter100|0931_ ;
  assign \new_Sorter100|1032_  = \new_Sorter100|0932_  & \new_Sorter100|0933_ ;
  assign \new_Sorter100|1033_  = \new_Sorter100|0932_  | \new_Sorter100|0933_ ;
  assign \new_Sorter100|1034_  = \new_Sorter100|0934_  & \new_Sorter100|0935_ ;
  assign \new_Sorter100|1035_  = \new_Sorter100|0934_  | \new_Sorter100|0935_ ;
  assign \new_Sorter100|1036_  = \new_Sorter100|0936_  & \new_Sorter100|0937_ ;
  assign \new_Sorter100|1037_  = \new_Sorter100|0936_  | \new_Sorter100|0937_ ;
  assign \new_Sorter100|1038_  = \new_Sorter100|0938_  & \new_Sorter100|0939_ ;
  assign \new_Sorter100|1039_  = \new_Sorter100|0938_  | \new_Sorter100|0939_ ;
  assign \new_Sorter100|1040_  = \new_Sorter100|0940_  & \new_Sorter100|0941_ ;
  assign \new_Sorter100|1041_  = \new_Sorter100|0940_  | \new_Sorter100|0941_ ;
  assign \new_Sorter100|1042_  = \new_Sorter100|0942_  & \new_Sorter100|0943_ ;
  assign \new_Sorter100|1043_  = \new_Sorter100|0942_  | \new_Sorter100|0943_ ;
  assign \new_Sorter100|1044_  = \new_Sorter100|0944_  & \new_Sorter100|0945_ ;
  assign \new_Sorter100|1045_  = \new_Sorter100|0944_  | \new_Sorter100|0945_ ;
  assign \new_Sorter100|1046_  = \new_Sorter100|0946_  & \new_Sorter100|0947_ ;
  assign \new_Sorter100|1047_  = \new_Sorter100|0946_  | \new_Sorter100|0947_ ;
  assign \new_Sorter100|1048_  = \new_Sorter100|0948_  & \new_Sorter100|0949_ ;
  assign \new_Sorter100|1049_  = \new_Sorter100|0948_  | \new_Sorter100|0949_ ;
  assign \new_Sorter100|1050_  = \new_Sorter100|0950_  & \new_Sorter100|0951_ ;
  assign \new_Sorter100|1051_  = \new_Sorter100|0950_  | \new_Sorter100|0951_ ;
  assign \new_Sorter100|1052_  = \new_Sorter100|0952_  & \new_Sorter100|0953_ ;
  assign \new_Sorter100|1053_  = \new_Sorter100|0952_  | \new_Sorter100|0953_ ;
  assign \new_Sorter100|1054_  = \new_Sorter100|0954_  & \new_Sorter100|0955_ ;
  assign \new_Sorter100|1055_  = \new_Sorter100|0954_  | \new_Sorter100|0955_ ;
  assign \new_Sorter100|1056_  = \new_Sorter100|0956_  & \new_Sorter100|0957_ ;
  assign \new_Sorter100|1057_  = \new_Sorter100|0956_  | \new_Sorter100|0957_ ;
  assign \new_Sorter100|1058_  = \new_Sorter100|0958_  & \new_Sorter100|0959_ ;
  assign \new_Sorter100|1059_  = \new_Sorter100|0958_  | \new_Sorter100|0959_ ;
  assign \new_Sorter100|1060_  = \new_Sorter100|0960_  & \new_Sorter100|0961_ ;
  assign \new_Sorter100|1061_  = \new_Sorter100|0960_  | \new_Sorter100|0961_ ;
  assign \new_Sorter100|1062_  = \new_Sorter100|0962_  & \new_Sorter100|0963_ ;
  assign \new_Sorter100|1063_  = \new_Sorter100|0962_  | \new_Sorter100|0963_ ;
  assign \new_Sorter100|1064_  = \new_Sorter100|0964_  & \new_Sorter100|0965_ ;
  assign \new_Sorter100|1065_  = \new_Sorter100|0964_  | \new_Sorter100|0965_ ;
  assign \new_Sorter100|1066_  = \new_Sorter100|0966_  & \new_Sorter100|0967_ ;
  assign \new_Sorter100|1067_  = \new_Sorter100|0966_  | \new_Sorter100|0967_ ;
  assign \new_Sorter100|1068_  = \new_Sorter100|0968_  & \new_Sorter100|0969_ ;
  assign \new_Sorter100|1069_  = \new_Sorter100|0968_  | \new_Sorter100|0969_ ;
  assign \new_Sorter100|1070_  = \new_Sorter100|0970_  & \new_Sorter100|0971_ ;
  assign \new_Sorter100|1071_  = \new_Sorter100|0970_  | \new_Sorter100|0971_ ;
  assign \new_Sorter100|1072_  = \new_Sorter100|0972_  & \new_Sorter100|0973_ ;
  assign \new_Sorter100|1073_  = \new_Sorter100|0972_  | \new_Sorter100|0973_ ;
  assign \new_Sorter100|1074_  = \new_Sorter100|0974_  & \new_Sorter100|0975_ ;
  assign \new_Sorter100|1075_  = \new_Sorter100|0974_  | \new_Sorter100|0975_ ;
  assign \new_Sorter100|1076_  = \new_Sorter100|0976_  & \new_Sorter100|0977_ ;
  assign \new_Sorter100|1077_  = \new_Sorter100|0976_  | \new_Sorter100|0977_ ;
  assign \new_Sorter100|1078_  = \new_Sorter100|0978_  & \new_Sorter100|0979_ ;
  assign \new_Sorter100|1079_  = \new_Sorter100|0978_  | \new_Sorter100|0979_ ;
  assign \new_Sorter100|1080_  = \new_Sorter100|0980_  & \new_Sorter100|0981_ ;
  assign \new_Sorter100|1081_  = \new_Sorter100|0980_  | \new_Sorter100|0981_ ;
  assign \new_Sorter100|1082_  = \new_Sorter100|0982_  & \new_Sorter100|0983_ ;
  assign \new_Sorter100|1083_  = \new_Sorter100|0982_  | \new_Sorter100|0983_ ;
  assign \new_Sorter100|1084_  = \new_Sorter100|0984_  & \new_Sorter100|0985_ ;
  assign \new_Sorter100|1085_  = \new_Sorter100|0984_  | \new_Sorter100|0985_ ;
  assign \new_Sorter100|1086_  = \new_Sorter100|0986_  & \new_Sorter100|0987_ ;
  assign \new_Sorter100|1087_  = \new_Sorter100|0986_  | \new_Sorter100|0987_ ;
  assign \new_Sorter100|1088_  = \new_Sorter100|0988_  & \new_Sorter100|0989_ ;
  assign \new_Sorter100|1089_  = \new_Sorter100|0988_  | \new_Sorter100|0989_ ;
  assign \new_Sorter100|1090_  = \new_Sorter100|0990_  & \new_Sorter100|0991_ ;
  assign \new_Sorter100|1091_  = \new_Sorter100|0990_  | \new_Sorter100|0991_ ;
  assign \new_Sorter100|1092_  = \new_Sorter100|0992_  & \new_Sorter100|0993_ ;
  assign \new_Sorter100|1093_  = \new_Sorter100|0992_  | \new_Sorter100|0993_ ;
  assign \new_Sorter100|1094_  = \new_Sorter100|0994_  & \new_Sorter100|0995_ ;
  assign \new_Sorter100|1095_  = \new_Sorter100|0994_  | \new_Sorter100|0995_ ;
  assign \new_Sorter100|1096_  = \new_Sorter100|0996_  & \new_Sorter100|0997_ ;
  assign \new_Sorter100|1097_  = \new_Sorter100|0996_  | \new_Sorter100|0997_ ;
  assign \new_Sorter100|1098_  = \new_Sorter100|0998_  & \new_Sorter100|0999_ ;
  assign \new_Sorter100|1099_  = \new_Sorter100|0998_  | \new_Sorter100|0999_ ;
  assign \new_Sorter100|1100_  = \new_Sorter100|1000_ ;
  assign \new_Sorter100|1199_  = \new_Sorter100|1099_ ;
  assign \new_Sorter100|1101_  = \new_Sorter100|1001_  & \new_Sorter100|1002_ ;
  assign \new_Sorter100|1102_  = \new_Sorter100|1001_  | \new_Sorter100|1002_ ;
  assign \new_Sorter100|1103_  = \new_Sorter100|1003_  & \new_Sorter100|1004_ ;
  assign \new_Sorter100|1104_  = \new_Sorter100|1003_  | \new_Sorter100|1004_ ;
  assign \new_Sorter100|1105_  = \new_Sorter100|1005_  & \new_Sorter100|1006_ ;
  assign \new_Sorter100|1106_  = \new_Sorter100|1005_  | \new_Sorter100|1006_ ;
  assign \new_Sorter100|1107_  = \new_Sorter100|1007_  & \new_Sorter100|1008_ ;
  assign \new_Sorter100|1108_  = \new_Sorter100|1007_  | \new_Sorter100|1008_ ;
  assign \new_Sorter100|1109_  = \new_Sorter100|1009_  & \new_Sorter100|1010_ ;
  assign \new_Sorter100|1110_  = \new_Sorter100|1009_  | \new_Sorter100|1010_ ;
  assign \new_Sorter100|1111_  = \new_Sorter100|1011_  & \new_Sorter100|1012_ ;
  assign \new_Sorter100|1112_  = \new_Sorter100|1011_  | \new_Sorter100|1012_ ;
  assign \new_Sorter100|1113_  = \new_Sorter100|1013_  & \new_Sorter100|1014_ ;
  assign \new_Sorter100|1114_  = \new_Sorter100|1013_  | \new_Sorter100|1014_ ;
  assign \new_Sorter100|1115_  = \new_Sorter100|1015_  & \new_Sorter100|1016_ ;
  assign \new_Sorter100|1116_  = \new_Sorter100|1015_  | \new_Sorter100|1016_ ;
  assign \new_Sorter100|1117_  = \new_Sorter100|1017_  & \new_Sorter100|1018_ ;
  assign \new_Sorter100|1118_  = \new_Sorter100|1017_  | \new_Sorter100|1018_ ;
  assign \new_Sorter100|1119_  = \new_Sorter100|1019_  & \new_Sorter100|1020_ ;
  assign \new_Sorter100|1120_  = \new_Sorter100|1019_  | \new_Sorter100|1020_ ;
  assign \new_Sorter100|1121_  = \new_Sorter100|1021_  & \new_Sorter100|1022_ ;
  assign \new_Sorter100|1122_  = \new_Sorter100|1021_  | \new_Sorter100|1022_ ;
  assign \new_Sorter100|1123_  = \new_Sorter100|1023_  & \new_Sorter100|1024_ ;
  assign \new_Sorter100|1124_  = \new_Sorter100|1023_  | \new_Sorter100|1024_ ;
  assign \new_Sorter100|1125_  = \new_Sorter100|1025_  & \new_Sorter100|1026_ ;
  assign \new_Sorter100|1126_  = \new_Sorter100|1025_  | \new_Sorter100|1026_ ;
  assign \new_Sorter100|1127_  = \new_Sorter100|1027_  & \new_Sorter100|1028_ ;
  assign \new_Sorter100|1128_  = \new_Sorter100|1027_  | \new_Sorter100|1028_ ;
  assign \new_Sorter100|1129_  = \new_Sorter100|1029_  & \new_Sorter100|1030_ ;
  assign \new_Sorter100|1130_  = \new_Sorter100|1029_  | \new_Sorter100|1030_ ;
  assign \new_Sorter100|1131_  = \new_Sorter100|1031_  & \new_Sorter100|1032_ ;
  assign \new_Sorter100|1132_  = \new_Sorter100|1031_  | \new_Sorter100|1032_ ;
  assign \new_Sorter100|1133_  = \new_Sorter100|1033_  & \new_Sorter100|1034_ ;
  assign \new_Sorter100|1134_  = \new_Sorter100|1033_  | \new_Sorter100|1034_ ;
  assign \new_Sorter100|1135_  = \new_Sorter100|1035_  & \new_Sorter100|1036_ ;
  assign \new_Sorter100|1136_  = \new_Sorter100|1035_  | \new_Sorter100|1036_ ;
  assign \new_Sorter100|1137_  = \new_Sorter100|1037_  & \new_Sorter100|1038_ ;
  assign \new_Sorter100|1138_  = \new_Sorter100|1037_  | \new_Sorter100|1038_ ;
  assign \new_Sorter100|1139_  = \new_Sorter100|1039_  & \new_Sorter100|1040_ ;
  assign \new_Sorter100|1140_  = \new_Sorter100|1039_  | \new_Sorter100|1040_ ;
  assign \new_Sorter100|1141_  = \new_Sorter100|1041_  & \new_Sorter100|1042_ ;
  assign \new_Sorter100|1142_  = \new_Sorter100|1041_  | \new_Sorter100|1042_ ;
  assign \new_Sorter100|1143_  = \new_Sorter100|1043_  & \new_Sorter100|1044_ ;
  assign \new_Sorter100|1144_  = \new_Sorter100|1043_  | \new_Sorter100|1044_ ;
  assign \new_Sorter100|1145_  = \new_Sorter100|1045_  & \new_Sorter100|1046_ ;
  assign \new_Sorter100|1146_  = \new_Sorter100|1045_  | \new_Sorter100|1046_ ;
  assign \new_Sorter100|1147_  = \new_Sorter100|1047_  & \new_Sorter100|1048_ ;
  assign \new_Sorter100|1148_  = \new_Sorter100|1047_  | \new_Sorter100|1048_ ;
  assign \new_Sorter100|1149_  = \new_Sorter100|1049_  & \new_Sorter100|1050_ ;
  assign \new_Sorter100|1150_  = \new_Sorter100|1049_  | \new_Sorter100|1050_ ;
  assign \new_Sorter100|1151_  = \new_Sorter100|1051_  & \new_Sorter100|1052_ ;
  assign \new_Sorter100|1152_  = \new_Sorter100|1051_  | \new_Sorter100|1052_ ;
  assign \new_Sorter100|1153_  = \new_Sorter100|1053_  & \new_Sorter100|1054_ ;
  assign \new_Sorter100|1154_  = \new_Sorter100|1053_  | \new_Sorter100|1054_ ;
  assign \new_Sorter100|1155_  = \new_Sorter100|1055_  & \new_Sorter100|1056_ ;
  assign \new_Sorter100|1156_  = \new_Sorter100|1055_  | \new_Sorter100|1056_ ;
  assign \new_Sorter100|1157_  = \new_Sorter100|1057_  & \new_Sorter100|1058_ ;
  assign \new_Sorter100|1158_  = \new_Sorter100|1057_  | \new_Sorter100|1058_ ;
  assign \new_Sorter100|1159_  = \new_Sorter100|1059_  & \new_Sorter100|1060_ ;
  assign \new_Sorter100|1160_  = \new_Sorter100|1059_  | \new_Sorter100|1060_ ;
  assign \new_Sorter100|1161_  = \new_Sorter100|1061_  & \new_Sorter100|1062_ ;
  assign \new_Sorter100|1162_  = \new_Sorter100|1061_  | \new_Sorter100|1062_ ;
  assign \new_Sorter100|1163_  = \new_Sorter100|1063_  & \new_Sorter100|1064_ ;
  assign \new_Sorter100|1164_  = \new_Sorter100|1063_  | \new_Sorter100|1064_ ;
  assign \new_Sorter100|1165_  = \new_Sorter100|1065_  & \new_Sorter100|1066_ ;
  assign \new_Sorter100|1166_  = \new_Sorter100|1065_  | \new_Sorter100|1066_ ;
  assign \new_Sorter100|1167_  = \new_Sorter100|1067_  & \new_Sorter100|1068_ ;
  assign \new_Sorter100|1168_  = \new_Sorter100|1067_  | \new_Sorter100|1068_ ;
  assign \new_Sorter100|1169_  = \new_Sorter100|1069_  & \new_Sorter100|1070_ ;
  assign \new_Sorter100|1170_  = \new_Sorter100|1069_  | \new_Sorter100|1070_ ;
  assign \new_Sorter100|1171_  = \new_Sorter100|1071_  & \new_Sorter100|1072_ ;
  assign \new_Sorter100|1172_  = \new_Sorter100|1071_  | \new_Sorter100|1072_ ;
  assign \new_Sorter100|1173_  = \new_Sorter100|1073_  & \new_Sorter100|1074_ ;
  assign \new_Sorter100|1174_  = \new_Sorter100|1073_  | \new_Sorter100|1074_ ;
  assign \new_Sorter100|1175_  = \new_Sorter100|1075_  & \new_Sorter100|1076_ ;
  assign \new_Sorter100|1176_  = \new_Sorter100|1075_  | \new_Sorter100|1076_ ;
  assign \new_Sorter100|1177_  = \new_Sorter100|1077_  & \new_Sorter100|1078_ ;
  assign \new_Sorter100|1178_  = \new_Sorter100|1077_  | \new_Sorter100|1078_ ;
  assign \new_Sorter100|1179_  = \new_Sorter100|1079_  & \new_Sorter100|1080_ ;
  assign \new_Sorter100|1180_  = \new_Sorter100|1079_  | \new_Sorter100|1080_ ;
  assign \new_Sorter100|1181_  = \new_Sorter100|1081_  & \new_Sorter100|1082_ ;
  assign \new_Sorter100|1182_  = \new_Sorter100|1081_  | \new_Sorter100|1082_ ;
  assign \new_Sorter100|1183_  = \new_Sorter100|1083_  & \new_Sorter100|1084_ ;
  assign \new_Sorter100|1184_  = \new_Sorter100|1083_  | \new_Sorter100|1084_ ;
  assign \new_Sorter100|1185_  = \new_Sorter100|1085_  & \new_Sorter100|1086_ ;
  assign \new_Sorter100|1186_  = \new_Sorter100|1085_  | \new_Sorter100|1086_ ;
  assign \new_Sorter100|1187_  = \new_Sorter100|1087_  & \new_Sorter100|1088_ ;
  assign \new_Sorter100|1188_  = \new_Sorter100|1087_  | \new_Sorter100|1088_ ;
  assign \new_Sorter100|1189_  = \new_Sorter100|1089_  & \new_Sorter100|1090_ ;
  assign \new_Sorter100|1190_  = \new_Sorter100|1089_  | \new_Sorter100|1090_ ;
  assign \new_Sorter100|1191_  = \new_Sorter100|1091_  & \new_Sorter100|1092_ ;
  assign \new_Sorter100|1192_  = \new_Sorter100|1091_  | \new_Sorter100|1092_ ;
  assign \new_Sorter100|1193_  = \new_Sorter100|1093_  & \new_Sorter100|1094_ ;
  assign \new_Sorter100|1194_  = \new_Sorter100|1093_  | \new_Sorter100|1094_ ;
  assign \new_Sorter100|1195_  = \new_Sorter100|1095_  & \new_Sorter100|1096_ ;
  assign \new_Sorter100|1196_  = \new_Sorter100|1095_  | \new_Sorter100|1096_ ;
  assign \new_Sorter100|1197_  = \new_Sorter100|1097_  & \new_Sorter100|1098_ ;
  assign \new_Sorter100|1198_  = \new_Sorter100|1097_  | \new_Sorter100|1098_ ;
  assign \new_Sorter100|1200_  = \new_Sorter100|1100_  & \new_Sorter100|1101_ ;
  assign \new_Sorter100|1201_  = \new_Sorter100|1100_  | \new_Sorter100|1101_ ;
  assign \new_Sorter100|1202_  = \new_Sorter100|1102_  & \new_Sorter100|1103_ ;
  assign \new_Sorter100|1203_  = \new_Sorter100|1102_  | \new_Sorter100|1103_ ;
  assign \new_Sorter100|1204_  = \new_Sorter100|1104_  & \new_Sorter100|1105_ ;
  assign \new_Sorter100|1205_  = \new_Sorter100|1104_  | \new_Sorter100|1105_ ;
  assign \new_Sorter100|1206_  = \new_Sorter100|1106_  & \new_Sorter100|1107_ ;
  assign \new_Sorter100|1207_  = \new_Sorter100|1106_  | \new_Sorter100|1107_ ;
  assign \new_Sorter100|1208_  = \new_Sorter100|1108_  & \new_Sorter100|1109_ ;
  assign \new_Sorter100|1209_  = \new_Sorter100|1108_  | \new_Sorter100|1109_ ;
  assign \new_Sorter100|1210_  = \new_Sorter100|1110_  & \new_Sorter100|1111_ ;
  assign \new_Sorter100|1211_  = \new_Sorter100|1110_  | \new_Sorter100|1111_ ;
  assign \new_Sorter100|1212_  = \new_Sorter100|1112_  & \new_Sorter100|1113_ ;
  assign \new_Sorter100|1213_  = \new_Sorter100|1112_  | \new_Sorter100|1113_ ;
  assign \new_Sorter100|1214_  = \new_Sorter100|1114_  & \new_Sorter100|1115_ ;
  assign \new_Sorter100|1215_  = \new_Sorter100|1114_  | \new_Sorter100|1115_ ;
  assign \new_Sorter100|1216_  = \new_Sorter100|1116_  & \new_Sorter100|1117_ ;
  assign \new_Sorter100|1217_  = \new_Sorter100|1116_  | \new_Sorter100|1117_ ;
  assign \new_Sorter100|1218_  = \new_Sorter100|1118_  & \new_Sorter100|1119_ ;
  assign \new_Sorter100|1219_  = \new_Sorter100|1118_  | \new_Sorter100|1119_ ;
  assign \new_Sorter100|1220_  = \new_Sorter100|1120_  & \new_Sorter100|1121_ ;
  assign \new_Sorter100|1221_  = \new_Sorter100|1120_  | \new_Sorter100|1121_ ;
  assign \new_Sorter100|1222_  = \new_Sorter100|1122_  & \new_Sorter100|1123_ ;
  assign \new_Sorter100|1223_  = \new_Sorter100|1122_  | \new_Sorter100|1123_ ;
  assign \new_Sorter100|1224_  = \new_Sorter100|1124_  & \new_Sorter100|1125_ ;
  assign \new_Sorter100|1225_  = \new_Sorter100|1124_  | \new_Sorter100|1125_ ;
  assign \new_Sorter100|1226_  = \new_Sorter100|1126_  & \new_Sorter100|1127_ ;
  assign \new_Sorter100|1227_  = \new_Sorter100|1126_  | \new_Sorter100|1127_ ;
  assign \new_Sorter100|1228_  = \new_Sorter100|1128_  & \new_Sorter100|1129_ ;
  assign \new_Sorter100|1229_  = \new_Sorter100|1128_  | \new_Sorter100|1129_ ;
  assign \new_Sorter100|1230_  = \new_Sorter100|1130_  & \new_Sorter100|1131_ ;
  assign \new_Sorter100|1231_  = \new_Sorter100|1130_  | \new_Sorter100|1131_ ;
  assign \new_Sorter100|1232_  = \new_Sorter100|1132_  & \new_Sorter100|1133_ ;
  assign \new_Sorter100|1233_  = \new_Sorter100|1132_  | \new_Sorter100|1133_ ;
  assign \new_Sorter100|1234_  = \new_Sorter100|1134_  & \new_Sorter100|1135_ ;
  assign \new_Sorter100|1235_  = \new_Sorter100|1134_  | \new_Sorter100|1135_ ;
  assign \new_Sorter100|1236_  = \new_Sorter100|1136_  & \new_Sorter100|1137_ ;
  assign \new_Sorter100|1237_  = \new_Sorter100|1136_  | \new_Sorter100|1137_ ;
  assign \new_Sorter100|1238_  = \new_Sorter100|1138_  & \new_Sorter100|1139_ ;
  assign \new_Sorter100|1239_  = \new_Sorter100|1138_  | \new_Sorter100|1139_ ;
  assign \new_Sorter100|1240_  = \new_Sorter100|1140_  & \new_Sorter100|1141_ ;
  assign \new_Sorter100|1241_  = \new_Sorter100|1140_  | \new_Sorter100|1141_ ;
  assign \new_Sorter100|1242_  = \new_Sorter100|1142_  & \new_Sorter100|1143_ ;
  assign \new_Sorter100|1243_  = \new_Sorter100|1142_  | \new_Sorter100|1143_ ;
  assign \new_Sorter100|1244_  = \new_Sorter100|1144_  & \new_Sorter100|1145_ ;
  assign \new_Sorter100|1245_  = \new_Sorter100|1144_  | \new_Sorter100|1145_ ;
  assign \new_Sorter100|1246_  = \new_Sorter100|1146_  & \new_Sorter100|1147_ ;
  assign \new_Sorter100|1247_  = \new_Sorter100|1146_  | \new_Sorter100|1147_ ;
  assign \new_Sorter100|1248_  = \new_Sorter100|1148_  & \new_Sorter100|1149_ ;
  assign \new_Sorter100|1249_  = \new_Sorter100|1148_  | \new_Sorter100|1149_ ;
  assign \new_Sorter100|1250_  = \new_Sorter100|1150_  & \new_Sorter100|1151_ ;
  assign \new_Sorter100|1251_  = \new_Sorter100|1150_  | \new_Sorter100|1151_ ;
  assign \new_Sorter100|1252_  = \new_Sorter100|1152_  & \new_Sorter100|1153_ ;
  assign \new_Sorter100|1253_  = \new_Sorter100|1152_  | \new_Sorter100|1153_ ;
  assign \new_Sorter100|1254_  = \new_Sorter100|1154_  & \new_Sorter100|1155_ ;
  assign \new_Sorter100|1255_  = \new_Sorter100|1154_  | \new_Sorter100|1155_ ;
  assign \new_Sorter100|1256_  = \new_Sorter100|1156_  & \new_Sorter100|1157_ ;
  assign \new_Sorter100|1257_  = \new_Sorter100|1156_  | \new_Sorter100|1157_ ;
  assign \new_Sorter100|1258_  = \new_Sorter100|1158_  & \new_Sorter100|1159_ ;
  assign \new_Sorter100|1259_  = \new_Sorter100|1158_  | \new_Sorter100|1159_ ;
  assign \new_Sorter100|1260_  = \new_Sorter100|1160_  & \new_Sorter100|1161_ ;
  assign \new_Sorter100|1261_  = \new_Sorter100|1160_  | \new_Sorter100|1161_ ;
  assign \new_Sorter100|1262_  = \new_Sorter100|1162_  & \new_Sorter100|1163_ ;
  assign \new_Sorter100|1263_  = \new_Sorter100|1162_  | \new_Sorter100|1163_ ;
  assign \new_Sorter100|1264_  = \new_Sorter100|1164_  & \new_Sorter100|1165_ ;
  assign \new_Sorter100|1265_  = \new_Sorter100|1164_  | \new_Sorter100|1165_ ;
  assign \new_Sorter100|1266_  = \new_Sorter100|1166_  & \new_Sorter100|1167_ ;
  assign \new_Sorter100|1267_  = \new_Sorter100|1166_  | \new_Sorter100|1167_ ;
  assign \new_Sorter100|1268_  = \new_Sorter100|1168_  & \new_Sorter100|1169_ ;
  assign \new_Sorter100|1269_  = \new_Sorter100|1168_  | \new_Sorter100|1169_ ;
  assign \new_Sorter100|1270_  = \new_Sorter100|1170_  & \new_Sorter100|1171_ ;
  assign \new_Sorter100|1271_  = \new_Sorter100|1170_  | \new_Sorter100|1171_ ;
  assign \new_Sorter100|1272_  = \new_Sorter100|1172_  & \new_Sorter100|1173_ ;
  assign \new_Sorter100|1273_  = \new_Sorter100|1172_  | \new_Sorter100|1173_ ;
  assign \new_Sorter100|1274_  = \new_Sorter100|1174_  & \new_Sorter100|1175_ ;
  assign \new_Sorter100|1275_  = \new_Sorter100|1174_  | \new_Sorter100|1175_ ;
  assign \new_Sorter100|1276_  = \new_Sorter100|1176_  & \new_Sorter100|1177_ ;
  assign \new_Sorter100|1277_  = \new_Sorter100|1176_  | \new_Sorter100|1177_ ;
  assign \new_Sorter100|1278_  = \new_Sorter100|1178_  & \new_Sorter100|1179_ ;
  assign \new_Sorter100|1279_  = \new_Sorter100|1178_  | \new_Sorter100|1179_ ;
  assign \new_Sorter100|1280_  = \new_Sorter100|1180_  & \new_Sorter100|1181_ ;
  assign \new_Sorter100|1281_  = \new_Sorter100|1180_  | \new_Sorter100|1181_ ;
  assign \new_Sorter100|1282_  = \new_Sorter100|1182_  & \new_Sorter100|1183_ ;
  assign \new_Sorter100|1283_  = \new_Sorter100|1182_  | \new_Sorter100|1183_ ;
  assign \new_Sorter100|1284_  = \new_Sorter100|1184_  & \new_Sorter100|1185_ ;
  assign \new_Sorter100|1285_  = \new_Sorter100|1184_  | \new_Sorter100|1185_ ;
  assign \new_Sorter100|1286_  = \new_Sorter100|1186_  & \new_Sorter100|1187_ ;
  assign \new_Sorter100|1287_  = \new_Sorter100|1186_  | \new_Sorter100|1187_ ;
  assign \new_Sorter100|1288_  = \new_Sorter100|1188_  & \new_Sorter100|1189_ ;
  assign \new_Sorter100|1289_  = \new_Sorter100|1188_  | \new_Sorter100|1189_ ;
  assign \new_Sorter100|1290_  = \new_Sorter100|1190_  & \new_Sorter100|1191_ ;
  assign \new_Sorter100|1291_  = \new_Sorter100|1190_  | \new_Sorter100|1191_ ;
  assign \new_Sorter100|1292_  = \new_Sorter100|1192_  & \new_Sorter100|1193_ ;
  assign \new_Sorter100|1293_  = \new_Sorter100|1192_  | \new_Sorter100|1193_ ;
  assign \new_Sorter100|1294_  = \new_Sorter100|1194_  & \new_Sorter100|1195_ ;
  assign \new_Sorter100|1295_  = \new_Sorter100|1194_  | \new_Sorter100|1195_ ;
  assign \new_Sorter100|1296_  = \new_Sorter100|1196_  & \new_Sorter100|1197_ ;
  assign \new_Sorter100|1297_  = \new_Sorter100|1196_  | \new_Sorter100|1197_ ;
  assign \new_Sorter100|1298_  = \new_Sorter100|1198_  & \new_Sorter100|1199_ ;
  assign \new_Sorter100|1299_  = \new_Sorter100|1198_  | \new_Sorter100|1199_ ;
  assign \new_Sorter100|1300_  = \new_Sorter100|1200_ ;
  assign \new_Sorter100|1399_  = \new_Sorter100|1299_ ;
  assign \new_Sorter100|1301_  = \new_Sorter100|1201_  & \new_Sorter100|1202_ ;
  assign \new_Sorter100|1302_  = \new_Sorter100|1201_  | \new_Sorter100|1202_ ;
  assign \new_Sorter100|1303_  = \new_Sorter100|1203_  & \new_Sorter100|1204_ ;
  assign \new_Sorter100|1304_  = \new_Sorter100|1203_  | \new_Sorter100|1204_ ;
  assign \new_Sorter100|1305_  = \new_Sorter100|1205_  & \new_Sorter100|1206_ ;
  assign \new_Sorter100|1306_  = \new_Sorter100|1205_  | \new_Sorter100|1206_ ;
  assign \new_Sorter100|1307_  = \new_Sorter100|1207_  & \new_Sorter100|1208_ ;
  assign \new_Sorter100|1308_  = \new_Sorter100|1207_  | \new_Sorter100|1208_ ;
  assign \new_Sorter100|1309_  = \new_Sorter100|1209_  & \new_Sorter100|1210_ ;
  assign \new_Sorter100|1310_  = \new_Sorter100|1209_  | \new_Sorter100|1210_ ;
  assign \new_Sorter100|1311_  = \new_Sorter100|1211_  & \new_Sorter100|1212_ ;
  assign \new_Sorter100|1312_  = \new_Sorter100|1211_  | \new_Sorter100|1212_ ;
  assign \new_Sorter100|1313_  = \new_Sorter100|1213_  & \new_Sorter100|1214_ ;
  assign \new_Sorter100|1314_  = \new_Sorter100|1213_  | \new_Sorter100|1214_ ;
  assign \new_Sorter100|1315_  = \new_Sorter100|1215_  & \new_Sorter100|1216_ ;
  assign \new_Sorter100|1316_  = \new_Sorter100|1215_  | \new_Sorter100|1216_ ;
  assign \new_Sorter100|1317_  = \new_Sorter100|1217_  & \new_Sorter100|1218_ ;
  assign \new_Sorter100|1318_  = \new_Sorter100|1217_  | \new_Sorter100|1218_ ;
  assign \new_Sorter100|1319_  = \new_Sorter100|1219_  & \new_Sorter100|1220_ ;
  assign \new_Sorter100|1320_  = \new_Sorter100|1219_  | \new_Sorter100|1220_ ;
  assign \new_Sorter100|1321_  = \new_Sorter100|1221_  & \new_Sorter100|1222_ ;
  assign \new_Sorter100|1322_  = \new_Sorter100|1221_  | \new_Sorter100|1222_ ;
  assign \new_Sorter100|1323_  = \new_Sorter100|1223_  & \new_Sorter100|1224_ ;
  assign \new_Sorter100|1324_  = \new_Sorter100|1223_  | \new_Sorter100|1224_ ;
  assign \new_Sorter100|1325_  = \new_Sorter100|1225_  & \new_Sorter100|1226_ ;
  assign \new_Sorter100|1326_  = \new_Sorter100|1225_  | \new_Sorter100|1226_ ;
  assign \new_Sorter100|1327_  = \new_Sorter100|1227_  & \new_Sorter100|1228_ ;
  assign \new_Sorter100|1328_  = \new_Sorter100|1227_  | \new_Sorter100|1228_ ;
  assign \new_Sorter100|1329_  = \new_Sorter100|1229_  & \new_Sorter100|1230_ ;
  assign \new_Sorter100|1330_  = \new_Sorter100|1229_  | \new_Sorter100|1230_ ;
  assign \new_Sorter100|1331_  = \new_Sorter100|1231_  & \new_Sorter100|1232_ ;
  assign \new_Sorter100|1332_  = \new_Sorter100|1231_  | \new_Sorter100|1232_ ;
  assign \new_Sorter100|1333_  = \new_Sorter100|1233_  & \new_Sorter100|1234_ ;
  assign \new_Sorter100|1334_  = \new_Sorter100|1233_  | \new_Sorter100|1234_ ;
  assign \new_Sorter100|1335_  = \new_Sorter100|1235_  & \new_Sorter100|1236_ ;
  assign \new_Sorter100|1336_  = \new_Sorter100|1235_  | \new_Sorter100|1236_ ;
  assign \new_Sorter100|1337_  = \new_Sorter100|1237_  & \new_Sorter100|1238_ ;
  assign \new_Sorter100|1338_  = \new_Sorter100|1237_  | \new_Sorter100|1238_ ;
  assign \new_Sorter100|1339_  = \new_Sorter100|1239_  & \new_Sorter100|1240_ ;
  assign \new_Sorter100|1340_  = \new_Sorter100|1239_  | \new_Sorter100|1240_ ;
  assign \new_Sorter100|1341_  = \new_Sorter100|1241_  & \new_Sorter100|1242_ ;
  assign \new_Sorter100|1342_  = \new_Sorter100|1241_  | \new_Sorter100|1242_ ;
  assign \new_Sorter100|1343_  = \new_Sorter100|1243_  & \new_Sorter100|1244_ ;
  assign \new_Sorter100|1344_  = \new_Sorter100|1243_  | \new_Sorter100|1244_ ;
  assign \new_Sorter100|1345_  = \new_Sorter100|1245_  & \new_Sorter100|1246_ ;
  assign \new_Sorter100|1346_  = \new_Sorter100|1245_  | \new_Sorter100|1246_ ;
  assign \new_Sorter100|1347_  = \new_Sorter100|1247_  & \new_Sorter100|1248_ ;
  assign \new_Sorter100|1348_  = \new_Sorter100|1247_  | \new_Sorter100|1248_ ;
  assign \new_Sorter100|1349_  = \new_Sorter100|1249_  & \new_Sorter100|1250_ ;
  assign \new_Sorter100|1350_  = \new_Sorter100|1249_  | \new_Sorter100|1250_ ;
  assign \new_Sorter100|1351_  = \new_Sorter100|1251_  & \new_Sorter100|1252_ ;
  assign \new_Sorter100|1352_  = \new_Sorter100|1251_  | \new_Sorter100|1252_ ;
  assign \new_Sorter100|1353_  = \new_Sorter100|1253_  & \new_Sorter100|1254_ ;
  assign \new_Sorter100|1354_  = \new_Sorter100|1253_  | \new_Sorter100|1254_ ;
  assign \new_Sorter100|1355_  = \new_Sorter100|1255_  & \new_Sorter100|1256_ ;
  assign \new_Sorter100|1356_  = \new_Sorter100|1255_  | \new_Sorter100|1256_ ;
  assign \new_Sorter100|1357_  = \new_Sorter100|1257_  & \new_Sorter100|1258_ ;
  assign \new_Sorter100|1358_  = \new_Sorter100|1257_  | \new_Sorter100|1258_ ;
  assign \new_Sorter100|1359_  = \new_Sorter100|1259_  & \new_Sorter100|1260_ ;
  assign \new_Sorter100|1360_  = \new_Sorter100|1259_  | \new_Sorter100|1260_ ;
  assign \new_Sorter100|1361_  = \new_Sorter100|1261_  & \new_Sorter100|1262_ ;
  assign \new_Sorter100|1362_  = \new_Sorter100|1261_  | \new_Sorter100|1262_ ;
  assign \new_Sorter100|1363_  = \new_Sorter100|1263_  & \new_Sorter100|1264_ ;
  assign \new_Sorter100|1364_  = \new_Sorter100|1263_  | \new_Sorter100|1264_ ;
  assign \new_Sorter100|1365_  = \new_Sorter100|1265_  & \new_Sorter100|1266_ ;
  assign \new_Sorter100|1366_  = \new_Sorter100|1265_  | \new_Sorter100|1266_ ;
  assign \new_Sorter100|1367_  = \new_Sorter100|1267_  & \new_Sorter100|1268_ ;
  assign \new_Sorter100|1368_  = \new_Sorter100|1267_  | \new_Sorter100|1268_ ;
  assign \new_Sorter100|1369_  = \new_Sorter100|1269_  & \new_Sorter100|1270_ ;
  assign \new_Sorter100|1370_  = \new_Sorter100|1269_  | \new_Sorter100|1270_ ;
  assign \new_Sorter100|1371_  = \new_Sorter100|1271_  & \new_Sorter100|1272_ ;
  assign \new_Sorter100|1372_  = \new_Sorter100|1271_  | \new_Sorter100|1272_ ;
  assign \new_Sorter100|1373_  = \new_Sorter100|1273_  & \new_Sorter100|1274_ ;
  assign \new_Sorter100|1374_  = \new_Sorter100|1273_  | \new_Sorter100|1274_ ;
  assign \new_Sorter100|1375_  = \new_Sorter100|1275_  & \new_Sorter100|1276_ ;
  assign \new_Sorter100|1376_  = \new_Sorter100|1275_  | \new_Sorter100|1276_ ;
  assign \new_Sorter100|1377_  = \new_Sorter100|1277_  & \new_Sorter100|1278_ ;
  assign \new_Sorter100|1378_  = \new_Sorter100|1277_  | \new_Sorter100|1278_ ;
  assign \new_Sorter100|1379_  = \new_Sorter100|1279_  & \new_Sorter100|1280_ ;
  assign \new_Sorter100|1380_  = \new_Sorter100|1279_  | \new_Sorter100|1280_ ;
  assign \new_Sorter100|1381_  = \new_Sorter100|1281_  & \new_Sorter100|1282_ ;
  assign \new_Sorter100|1382_  = \new_Sorter100|1281_  | \new_Sorter100|1282_ ;
  assign \new_Sorter100|1383_  = \new_Sorter100|1283_  & \new_Sorter100|1284_ ;
  assign \new_Sorter100|1384_  = \new_Sorter100|1283_  | \new_Sorter100|1284_ ;
  assign \new_Sorter100|1385_  = \new_Sorter100|1285_  & \new_Sorter100|1286_ ;
  assign \new_Sorter100|1386_  = \new_Sorter100|1285_  | \new_Sorter100|1286_ ;
  assign \new_Sorter100|1387_  = \new_Sorter100|1287_  & \new_Sorter100|1288_ ;
  assign \new_Sorter100|1388_  = \new_Sorter100|1287_  | \new_Sorter100|1288_ ;
  assign \new_Sorter100|1389_  = \new_Sorter100|1289_  & \new_Sorter100|1290_ ;
  assign \new_Sorter100|1390_  = \new_Sorter100|1289_  | \new_Sorter100|1290_ ;
  assign \new_Sorter100|1391_  = \new_Sorter100|1291_  & \new_Sorter100|1292_ ;
  assign \new_Sorter100|1392_  = \new_Sorter100|1291_  | \new_Sorter100|1292_ ;
  assign \new_Sorter100|1393_  = \new_Sorter100|1293_  & \new_Sorter100|1294_ ;
  assign \new_Sorter100|1394_  = \new_Sorter100|1293_  | \new_Sorter100|1294_ ;
  assign \new_Sorter100|1395_  = \new_Sorter100|1295_  & \new_Sorter100|1296_ ;
  assign \new_Sorter100|1396_  = \new_Sorter100|1295_  | \new_Sorter100|1296_ ;
  assign \new_Sorter100|1397_  = \new_Sorter100|1297_  & \new_Sorter100|1298_ ;
  assign \new_Sorter100|1398_  = \new_Sorter100|1297_  | \new_Sorter100|1298_ ;
  assign \new_Sorter100|1400_  = \new_Sorter100|1300_  & \new_Sorter100|1301_ ;
  assign \new_Sorter100|1401_  = \new_Sorter100|1300_  | \new_Sorter100|1301_ ;
  assign \new_Sorter100|1402_  = \new_Sorter100|1302_  & \new_Sorter100|1303_ ;
  assign \new_Sorter100|1403_  = \new_Sorter100|1302_  | \new_Sorter100|1303_ ;
  assign \new_Sorter100|1404_  = \new_Sorter100|1304_  & \new_Sorter100|1305_ ;
  assign \new_Sorter100|1405_  = \new_Sorter100|1304_  | \new_Sorter100|1305_ ;
  assign \new_Sorter100|1406_  = \new_Sorter100|1306_  & \new_Sorter100|1307_ ;
  assign \new_Sorter100|1407_  = \new_Sorter100|1306_  | \new_Sorter100|1307_ ;
  assign \new_Sorter100|1408_  = \new_Sorter100|1308_  & \new_Sorter100|1309_ ;
  assign \new_Sorter100|1409_  = \new_Sorter100|1308_  | \new_Sorter100|1309_ ;
  assign \new_Sorter100|1410_  = \new_Sorter100|1310_  & \new_Sorter100|1311_ ;
  assign \new_Sorter100|1411_  = \new_Sorter100|1310_  | \new_Sorter100|1311_ ;
  assign \new_Sorter100|1412_  = \new_Sorter100|1312_  & \new_Sorter100|1313_ ;
  assign \new_Sorter100|1413_  = \new_Sorter100|1312_  | \new_Sorter100|1313_ ;
  assign \new_Sorter100|1414_  = \new_Sorter100|1314_  & \new_Sorter100|1315_ ;
  assign \new_Sorter100|1415_  = \new_Sorter100|1314_  | \new_Sorter100|1315_ ;
  assign \new_Sorter100|1416_  = \new_Sorter100|1316_  & \new_Sorter100|1317_ ;
  assign \new_Sorter100|1417_  = \new_Sorter100|1316_  | \new_Sorter100|1317_ ;
  assign \new_Sorter100|1418_  = \new_Sorter100|1318_  & \new_Sorter100|1319_ ;
  assign \new_Sorter100|1419_  = \new_Sorter100|1318_  | \new_Sorter100|1319_ ;
  assign \new_Sorter100|1420_  = \new_Sorter100|1320_  & \new_Sorter100|1321_ ;
  assign \new_Sorter100|1421_  = \new_Sorter100|1320_  | \new_Sorter100|1321_ ;
  assign \new_Sorter100|1422_  = \new_Sorter100|1322_  & \new_Sorter100|1323_ ;
  assign \new_Sorter100|1423_  = \new_Sorter100|1322_  | \new_Sorter100|1323_ ;
  assign \new_Sorter100|1424_  = \new_Sorter100|1324_  & \new_Sorter100|1325_ ;
  assign \new_Sorter100|1425_  = \new_Sorter100|1324_  | \new_Sorter100|1325_ ;
  assign \new_Sorter100|1426_  = \new_Sorter100|1326_  & \new_Sorter100|1327_ ;
  assign \new_Sorter100|1427_  = \new_Sorter100|1326_  | \new_Sorter100|1327_ ;
  assign \new_Sorter100|1428_  = \new_Sorter100|1328_  & \new_Sorter100|1329_ ;
  assign \new_Sorter100|1429_  = \new_Sorter100|1328_  | \new_Sorter100|1329_ ;
  assign \new_Sorter100|1430_  = \new_Sorter100|1330_  & \new_Sorter100|1331_ ;
  assign \new_Sorter100|1431_  = \new_Sorter100|1330_  | \new_Sorter100|1331_ ;
  assign \new_Sorter100|1432_  = \new_Sorter100|1332_  & \new_Sorter100|1333_ ;
  assign \new_Sorter100|1433_  = \new_Sorter100|1332_  | \new_Sorter100|1333_ ;
  assign \new_Sorter100|1434_  = \new_Sorter100|1334_  & \new_Sorter100|1335_ ;
  assign \new_Sorter100|1435_  = \new_Sorter100|1334_  | \new_Sorter100|1335_ ;
  assign \new_Sorter100|1436_  = \new_Sorter100|1336_  & \new_Sorter100|1337_ ;
  assign \new_Sorter100|1437_  = \new_Sorter100|1336_  | \new_Sorter100|1337_ ;
  assign \new_Sorter100|1438_  = \new_Sorter100|1338_  & \new_Sorter100|1339_ ;
  assign \new_Sorter100|1439_  = \new_Sorter100|1338_  | \new_Sorter100|1339_ ;
  assign \new_Sorter100|1440_  = \new_Sorter100|1340_  & \new_Sorter100|1341_ ;
  assign \new_Sorter100|1441_  = \new_Sorter100|1340_  | \new_Sorter100|1341_ ;
  assign \new_Sorter100|1442_  = \new_Sorter100|1342_  & \new_Sorter100|1343_ ;
  assign \new_Sorter100|1443_  = \new_Sorter100|1342_  | \new_Sorter100|1343_ ;
  assign \new_Sorter100|1444_  = \new_Sorter100|1344_  & \new_Sorter100|1345_ ;
  assign \new_Sorter100|1445_  = \new_Sorter100|1344_  | \new_Sorter100|1345_ ;
  assign \new_Sorter100|1446_  = \new_Sorter100|1346_  & \new_Sorter100|1347_ ;
  assign \new_Sorter100|1447_  = \new_Sorter100|1346_  | \new_Sorter100|1347_ ;
  assign \new_Sorter100|1448_  = \new_Sorter100|1348_  & \new_Sorter100|1349_ ;
  assign \new_Sorter100|1449_  = \new_Sorter100|1348_  | \new_Sorter100|1349_ ;
  assign \new_Sorter100|1450_  = \new_Sorter100|1350_  & \new_Sorter100|1351_ ;
  assign \new_Sorter100|1451_  = \new_Sorter100|1350_  | \new_Sorter100|1351_ ;
  assign \new_Sorter100|1452_  = \new_Sorter100|1352_  & \new_Sorter100|1353_ ;
  assign \new_Sorter100|1453_  = \new_Sorter100|1352_  | \new_Sorter100|1353_ ;
  assign \new_Sorter100|1454_  = \new_Sorter100|1354_  & \new_Sorter100|1355_ ;
  assign \new_Sorter100|1455_  = \new_Sorter100|1354_  | \new_Sorter100|1355_ ;
  assign \new_Sorter100|1456_  = \new_Sorter100|1356_  & \new_Sorter100|1357_ ;
  assign \new_Sorter100|1457_  = \new_Sorter100|1356_  | \new_Sorter100|1357_ ;
  assign \new_Sorter100|1458_  = \new_Sorter100|1358_  & \new_Sorter100|1359_ ;
  assign \new_Sorter100|1459_  = \new_Sorter100|1358_  | \new_Sorter100|1359_ ;
  assign \new_Sorter100|1460_  = \new_Sorter100|1360_  & \new_Sorter100|1361_ ;
  assign \new_Sorter100|1461_  = \new_Sorter100|1360_  | \new_Sorter100|1361_ ;
  assign \new_Sorter100|1462_  = \new_Sorter100|1362_  & \new_Sorter100|1363_ ;
  assign \new_Sorter100|1463_  = \new_Sorter100|1362_  | \new_Sorter100|1363_ ;
  assign \new_Sorter100|1464_  = \new_Sorter100|1364_  & \new_Sorter100|1365_ ;
  assign \new_Sorter100|1465_  = \new_Sorter100|1364_  | \new_Sorter100|1365_ ;
  assign \new_Sorter100|1466_  = \new_Sorter100|1366_  & \new_Sorter100|1367_ ;
  assign \new_Sorter100|1467_  = \new_Sorter100|1366_  | \new_Sorter100|1367_ ;
  assign \new_Sorter100|1468_  = \new_Sorter100|1368_  & \new_Sorter100|1369_ ;
  assign \new_Sorter100|1469_  = \new_Sorter100|1368_  | \new_Sorter100|1369_ ;
  assign \new_Sorter100|1470_  = \new_Sorter100|1370_  & \new_Sorter100|1371_ ;
  assign \new_Sorter100|1471_  = \new_Sorter100|1370_  | \new_Sorter100|1371_ ;
  assign \new_Sorter100|1472_  = \new_Sorter100|1372_  & \new_Sorter100|1373_ ;
  assign \new_Sorter100|1473_  = \new_Sorter100|1372_  | \new_Sorter100|1373_ ;
  assign \new_Sorter100|1474_  = \new_Sorter100|1374_  & \new_Sorter100|1375_ ;
  assign \new_Sorter100|1475_  = \new_Sorter100|1374_  | \new_Sorter100|1375_ ;
  assign \new_Sorter100|1476_  = \new_Sorter100|1376_  & \new_Sorter100|1377_ ;
  assign \new_Sorter100|1477_  = \new_Sorter100|1376_  | \new_Sorter100|1377_ ;
  assign \new_Sorter100|1478_  = \new_Sorter100|1378_  & \new_Sorter100|1379_ ;
  assign \new_Sorter100|1479_  = \new_Sorter100|1378_  | \new_Sorter100|1379_ ;
  assign \new_Sorter100|1480_  = \new_Sorter100|1380_  & \new_Sorter100|1381_ ;
  assign \new_Sorter100|1481_  = \new_Sorter100|1380_  | \new_Sorter100|1381_ ;
  assign \new_Sorter100|1482_  = \new_Sorter100|1382_  & \new_Sorter100|1383_ ;
  assign \new_Sorter100|1483_  = \new_Sorter100|1382_  | \new_Sorter100|1383_ ;
  assign \new_Sorter100|1484_  = \new_Sorter100|1384_  & \new_Sorter100|1385_ ;
  assign \new_Sorter100|1485_  = \new_Sorter100|1384_  | \new_Sorter100|1385_ ;
  assign \new_Sorter100|1486_  = \new_Sorter100|1386_  & \new_Sorter100|1387_ ;
  assign \new_Sorter100|1487_  = \new_Sorter100|1386_  | \new_Sorter100|1387_ ;
  assign \new_Sorter100|1488_  = \new_Sorter100|1388_  & \new_Sorter100|1389_ ;
  assign \new_Sorter100|1489_  = \new_Sorter100|1388_  | \new_Sorter100|1389_ ;
  assign \new_Sorter100|1490_  = \new_Sorter100|1390_  & \new_Sorter100|1391_ ;
  assign \new_Sorter100|1491_  = \new_Sorter100|1390_  | \new_Sorter100|1391_ ;
  assign \new_Sorter100|1492_  = \new_Sorter100|1392_  & \new_Sorter100|1393_ ;
  assign \new_Sorter100|1493_  = \new_Sorter100|1392_  | \new_Sorter100|1393_ ;
  assign \new_Sorter100|1494_  = \new_Sorter100|1394_  & \new_Sorter100|1395_ ;
  assign \new_Sorter100|1495_  = \new_Sorter100|1394_  | \new_Sorter100|1395_ ;
  assign \new_Sorter100|1496_  = \new_Sorter100|1396_  & \new_Sorter100|1397_ ;
  assign \new_Sorter100|1497_  = \new_Sorter100|1396_  | \new_Sorter100|1397_ ;
  assign \new_Sorter100|1498_  = \new_Sorter100|1398_  & \new_Sorter100|1399_ ;
  assign \new_Sorter100|1499_  = \new_Sorter100|1398_  | \new_Sorter100|1399_ ;
  assign \new_Sorter100|1500_  = \new_Sorter100|1400_ ;
  assign \new_Sorter100|1599_  = \new_Sorter100|1499_ ;
  assign \new_Sorter100|1501_  = \new_Sorter100|1401_  & \new_Sorter100|1402_ ;
  assign \new_Sorter100|1502_  = \new_Sorter100|1401_  | \new_Sorter100|1402_ ;
  assign \new_Sorter100|1503_  = \new_Sorter100|1403_  & \new_Sorter100|1404_ ;
  assign \new_Sorter100|1504_  = \new_Sorter100|1403_  | \new_Sorter100|1404_ ;
  assign \new_Sorter100|1505_  = \new_Sorter100|1405_  & \new_Sorter100|1406_ ;
  assign \new_Sorter100|1506_  = \new_Sorter100|1405_  | \new_Sorter100|1406_ ;
  assign \new_Sorter100|1507_  = \new_Sorter100|1407_  & \new_Sorter100|1408_ ;
  assign \new_Sorter100|1508_  = \new_Sorter100|1407_  | \new_Sorter100|1408_ ;
  assign \new_Sorter100|1509_  = \new_Sorter100|1409_  & \new_Sorter100|1410_ ;
  assign \new_Sorter100|1510_  = \new_Sorter100|1409_  | \new_Sorter100|1410_ ;
  assign \new_Sorter100|1511_  = \new_Sorter100|1411_  & \new_Sorter100|1412_ ;
  assign \new_Sorter100|1512_  = \new_Sorter100|1411_  | \new_Sorter100|1412_ ;
  assign \new_Sorter100|1513_  = \new_Sorter100|1413_  & \new_Sorter100|1414_ ;
  assign \new_Sorter100|1514_  = \new_Sorter100|1413_  | \new_Sorter100|1414_ ;
  assign \new_Sorter100|1515_  = \new_Sorter100|1415_  & \new_Sorter100|1416_ ;
  assign \new_Sorter100|1516_  = \new_Sorter100|1415_  | \new_Sorter100|1416_ ;
  assign \new_Sorter100|1517_  = \new_Sorter100|1417_  & \new_Sorter100|1418_ ;
  assign \new_Sorter100|1518_  = \new_Sorter100|1417_  | \new_Sorter100|1418_ ;
  assign \new_Sorter100|1519_  = \new_Sorter100|1419_  & \new_Sorter100|1420_ ;
  assign \new_Sorter100|1520_  = \new_Sorter100|1419_  | \new_Sorter100|1420_ ;
  assign \new_Sorter100|1521_  = \new_Sorter100|1421_  & \new_Sorter100|1422_ ;
  assign \new_Sorter100|1522_  = \new_Sorter100|1421_  | \new_Sorter100|1422_ ;
  assign \new_Sorter100|1523_  = \new_Sorter100|1423_  & \new_Sorter100|1424_ ;
  assign \new_Sorter100|1524_  = \new_Sorter100|1423_  | \new_Sorter100|1424_ ;
  assign \new_Sorter100|1525_  = \new_Sorter100|1425_  & \new_Sorter100|1426_ ;
  assign \new_Sorter100|1526_  = \new_Sorter100|1425_  | \new_Sorter100|1426_ ;
  assign \new_Sorter100|1527_  = \new_Sorter100|1427_  & \new_Sorter100|1428_ ;
  assign \new_Sorter100|1528_  = \new_Sorter100|1427_  | \new_Sorter100|1428_ ;
  assign \new_Sorter100|1529_  = \new_Sorter100|1429_  & \new_Sorter100|1430_ ;
  assign \new_Sorter100|1530_  = \new_Sorter100|1429_  | \new_Sorter100|1430_ ;
  assign \new_Sorter100|1531_  = \new_Sorter100|1431_  & \new_Sorter100|1432_ ;
  assign \new_Sorter100|1532_  = \new_Sorter100|1431_  | \new_Sorter100|1432_ ;
  assign \new_Sorter100|1533_  = \new_Sorter100|1433_  & \new_Sorter100|1434_ ;
  assign \new_Sorter100|1534_  = \new_Sorter100|1433_  | \new_Sorter100|1434_ ;
  assign \new_Sorter100|1535_  = \new_Sorter100|1435_  & \new_Sorter100|1436_ ;
  assign \new_Sorter100|1536_  = \new_Sorter100|1435_  | \new_Sorter100|1436_ ;
  assign \new_Sorter100|1537_  = \new_Sorter100|1437_  & \new_Sorter100|1438_ ;
  assign \new_Sorter100|1538_  = \new_Sorter100|1437_  | \new_Sorter100|1438_ ;
  assign \new_Sorter100|1539_  = \new_Sorter100|1439_  & \new_Sorter100|1440_ ;
  assign \new_Sorter100|1540_  = \new_Sorter100|1439_  | \new_Sorter100|1440_ ;
  assign \new_Sorter100|1541_  = \new_Sorter100|1441_  & \new_Sorter100|1442_ ;
  assign \new_Sorter100|1542_  = \new_Sorter100|1441_  | \new_Sorter100|1442_ ;
  assign \new_Sorter100|1543_  = \new_Sorter100|1443_  & \new_Sorter100|1444_ ;
  assign \new_Sorter100|1544_  = \new_Sorter100|1443_  | \new_Sorter100|1444_ ;
  assign \new_Sorter100|1545_  = \new_Sorter100|1445_  & \new_Sorter100|1446_ ;
  assign \new_Sorter100|1546_  = \new_Sorter100|1445_  | \new_Sorter100|1446_ ;
  assign \new_Sorter100|1547_  = \new_Sorter100|1447_  & \new_Sorter100|1448_ ;
  assign \new_Sorter100|1548_  = \new_Sorter100|1447_  | \new_Sorter100|1448_ ;
  assign \new_Sorter100|1549_  = \new_Sorter100|1449_  & \new_Sorter100|1450_ ;
  assign \new_Sorter100|1550_  = \new_Sorter100|1449_  | \new_Sorter100|1450_ ;
  assign \new_Sorter100|1551_  = \new_Sorter100|1451_  & \new_Sorter100|1452_ ;
  assign \new_Sorter100|1552_  = \new_Sorter100|1451_  | \new_Sorter100|1452_ ;
  assign \new_Sorter100|1553_  = \new_Sorter100|1453_  & \new_Sorter100|1454_ ;
  assign \new_Sorter100|1554_  = \new_Sorter100|1453_  | \new_Sorter100|1454_ ;
  assign \new_Sorter100|1555_  = \new_Sorter100|1455_  & \new_Sorter100|1456_ ;
  assign \new_Sorter100|1556_  = \new_Sorter100|1455_  | \new_Sorter100|1456_ ;
  assign \new_Sorter100|1557_  = \new_Sorter100|1457_  & \new_Sorter100|1458_ ;
  assign \new_Sorter100|1558_  = \new_Sorter100|1457_  | \new_Sorter100|1458_ ;
  assign \new_Sorter100|1559_  = \new_Sorter100|1459_  & \new_Sorter100|1460_ ;
  assign \new_Sorter100|1560_  = \new_Sorter100|1459_  | \new_Sorter100|1460_ ;
  assign \new_Sorter100|1561_  = \new_Sorter100|1461_  & \new_Sorter100|1462_ ;
  assign \new_Sorter100|1562_  = \new_Sorter100|1461_  | \new_Sorter100|1462_ ;
  assign \new_Sorter100|1563_  = \new_Sorter100|1463_  & \new_Sorter100|1464_ ;
  assign \new_Sorter100|1564_  = \new_Sorter100|1463_  | \new_Sorter100|1464_ ;
  assign \new_Sorter100|1565_  = \new_Sorter100|1465_  & \new_Sorter100|1466_ ;
  assign \new_Sorter100|1566_  = \new_Sorter100|1465_  | \new_Sorter100|1466_ ;
  assign \new_Sorter100|1567_  = \new_Sorter100|1467_  & \new_Sorter100|1468_ ;
  assign \new_Sorter100|1568_  = \new_Sorter100|1467_  | \new_Sorter100|1468_ ;
  assign \new_Sorter100|1569_  = \new_Sorter100|1469_  & \new_Sorter100|1470_ ;
  assign \new_Sorter100|1570_  = \new_Sorter100|1469_  | \new_Sorter100|1470_ ;
  assign \new_Sorter100|1571_  = \new_Sorter100|1471_  & \new_Sorter100|1472_ ;
  assign \new_Sorter100|1572_  = \new_Sorter100|1471_  | \new_Sorter100|1472_ ;
  assign \new_Sorter100|1573_  = \new_Sorter100|1473_  & \new_Sorter100|1474_ ;
  assign \new_Sorter100|1574_  = \new_Sorter100|1473_  | \new_Sorter100|1474_ ;
  assign \new_Sorter100|1575_  = \new_Sorter100|1475_  & \new_Sorter100|1476_ ;
  assign \new_Sorter100|1576_  = \new_Sorter100|1475_  | \new_Sorter100|1476_ ;
  assign \new_Sorter100|1577_  = \new_Sorter100|1477_  & \new_Sorter100|1478_ ;
  assign \new_Sorter100|1578_  = \new_Sorter100|1477_  | \new_Sorter100|1478_ ;
  assign \new_Sorter100|1579_  = \new_Sorter100|1479_  & \new_Sorter100|1480_ ;
  assign \new_Sorter100|1580_  = \new_Sorter100|1479_  | \new_Sorter100|1480_ ;
  assign \new_Sorter100|1581_  = \new_Sorter100|1481_  & \new_Sorter100|1482_ ;
  assign \new_Sorter100|1582_  = \new_Sorter100|1481_  | \new_Sorter100|1482_ ;
  assign \new_Sorter100|1583_  = \new_Sorter100|1483_  & \new_Sorter100|1484_ ;
  assign \new_Sorter100|1584_  = \new_Sorter100|1483_  | \new_Sorter100|1484_ ;
  assign \new_Sorter100|1585_  = \new_Sorter100|1485_  & \new_Sorter100|1486_ ;
  assign \new_Sorter100|1586_  = \new_Sorter100|1485_  | \new_Sorter100|1486_ ;
  assign \new_Sorter100|1587_  = \new_Sorter100|1487_  & \new_Sorter100|1488_ ;
  assign \new_Sorter100|1588_  = \new_Sorter100|1487_  | \new_Sorter100|1488_ ;
  assign \new_Sorter100|1589_  = \new_Sorter100|1489_  & \new_Sorter100|1490_ ;
  assign \new_Sorter100|1590_  = \new_Sorter100|1489_  | \new_Sorter100|1490_ ;
  assign \new_Sorter100|1591_  = \new_Sorter100|1491_  & \new_Sorter100|1492_ ;
  assign \new_Sorter100|1592_  = \new_Sorter100|1491_  | \new_Sorter100|1492_ ;
  assign \new_Sorter100|1593_  = \new_Sorter100|1493_  & \new_Sorter100|1494_ ;
  assign \new_Sorter100|1594_  = \new_Sorter100|1493_  | \new_Sorter100|1494_ ;
  assign \new_Sorter100|1595_  = \new_Sorter100|1495_  & \new_Sorter100|1496_ ;
  assign \new_Sorter100|1596_  = \new_Sorter100|1495_  | \new_Sorter100|1496_ ;
  assign \new_Sorter100|1597_  = \new_Sorter100|1497_  & \new_Sorter100|1498_ ;
  assign \new_Sorter100|1598_  = \new_Sorter100|1497_  | \new_Sorter100|1498_ ;
  assign \new_Sorter100|1600_  = \new_Sorter100|1500_  & \new_Sorter100|1501_ ;
  assign \new_Sorter100|1601_  = \new_Sorter100|1500_  | \new_Sorter100|1501_ ;
  assign \new_Sorter100|1602_  = \new_Sorter100|1502_  & \new_Sorter100|1503_ ;
  assign \new_Sorter100|1603_  = \new_Sorter100|1502_  | \new_Sorter100|1503_ ;
  assign \new_Sorter100|1604_  = \new_Sorter100|1504_  & \new_Sorter100|1505_ ;
  assign \new_Sorter100|1605_  = \new_Sorter100|1504_  | \new_Sorter100|1505_ ;
  assign \new_Sorter100|1606_  = \new_Sorter100|1506_  & \new_Sorter100|1507_ ;
  assign \new_Sorter100|1607_  = \new_Sorter100|1506_  | \new_Sorter100|1507_ ;
  assign \new_Sorter100|1608_  = \new_Sorter100|1508_  & \new_Sorter100|1509_ ;
  assign \new_Sorter100|1609_  = \new_Sorter100|1508_  | \new_Sorter100|1509_ ;
  assign \new_Sorter100|1610_  = \new_Sorter100|1510_  & \new_Sorter100|1511_ ;
  assign \new_Sorter100|1611_  = \new_Sorter100|1510_  | \new_Sorter100|1511_ ;
  assign \new_Sorter100|1612_  = \new_Sorter100|1512_  & \new_Sorter100|1513_ ;
  assign \new_Sorter100|1613_  = \new_Sorter100|1512_  | \new_Sorter100|1513_ ;
  assign \new_Sorter100|1614_  = \new_Sorter100|1514_  & \new_Sorter100|1515_ ;
  assign \new_Sorter100|1615_  = \new_Sorter100|1514_  | \new_Sorter100|1515_ ;
  assign \new_Sorter100|1616_  = \new_Sorter100|1516_  & \new_Sorter100|1517_ ;
  assign \new_Sorter100|1617_  = \new_Sorter100|1516_  | \new_Sorter100|1517_ ;
  assign \new_Sorter100|1618_  = \new_Sorter100|1518_  & \new_Sorter100|1519_ ;
  assign \new_Sorter100|1619_  = \new_Sorter100|1518_  | \new_Sorter100|1519_ ;
  assign \new_Sorter100|1620_  = \new_Sorter100|1520_  & \new_Sorter100|1521_ ;
  assign \new_Sorter100|1621_  = \new_Sorter100|1520_  | \new_Sorter100|1521_ ;
  assign \new_Sorter100|1622_  = \new_Sorter100|1522_  & \new_Sorter100|1523_ ;
  assign \new_Sorter100|1623_  = \new_Sorter100|1522_  | \new_Sorter100|1523_ ;
  assign \new_Sorter100|1624_  = \new_Sorter100|1524_  & \new_Sorter100|1525_ ;
  assign \new_Sorter100|1625_  = \new_Sorter100|1524_  | \new_Sorter100|1525_ ;
  assign \new_Sorter100|1626_  = \new_Sorter100|1526_  & \new_Sorter100|1527_ ;
  assign \new_Sorter100|1627_  = \new_Sorter100|1526_  | \new_Sorter100|1527_ ;
  assign \new_Sorter100|1628_  = \new_Sorter100|1528_  & \new_Sorter100|1529_ ;
  assign \new_Sorter100|1629_  = \new_Sorter100|1528_  | \new_Sorter100|1529_ ;
  assign \new_Sorter100|1630_  = \new_Sorter100|1530_  & \new_Sorter100|1531_ ;
  assign \new_Sorter100|1631_  = \new_Sorter100|1530_  | \new_Sorter100|1531_ ;
  assign \new_Sorter100|1632_  = \new_Sorter100|1532_  & \new_Sorter100|1533_ ;
  assign \new_Sorter100|1633_  = \new_Sorter100|1532_  | \new_Sorter100|1533_ ;
  assign \new_Sorter100|1634_  = \new_Sorter100|1534_  & \new_Sorter100|1535_ ;
  assign \new_Sorter100|1635_  = \new_Sorter100|1534_  | \new_Sorter100|1535_ ;
  assign \new_Sorter100|1636_  = \new_Sorter100|1536_  & \new_Sorter100|1537_ ;
  assign \new_Sorter100|1637_  = \new_Sorter100|1536_  | \new_Sorter100|1537_ ;
  assign \new_Sorter100|1638_  = \new_Sorter100|1538_  & \new_Sorter100|1539_ ;
  assign \new_Sorter100|1639_  = \new_Sorter100|1538_  | \new_Sorter100|1539_ ;
  assign \new_Sorter100|1640_  = \new_Sorter100|1540_  & \new_Sorter100|1541_ ;
  assign \new_Sorter100|1641_  = \new_Sorter100|1540_  | \new_Sorter100|1541_ ;
  assign \new_Sorter100|1642_  = \new_Sorter100|1542_  & \new_Sorter100|1543_ ;
  assign \new_Sorter100|1643_  = \new_Sorter100|1542_  | \new_Sorter100|1543_ ;
  assign \new_Sorter100|1644_  = \new_Sorter100|1544_  & \new_Sorter100|1545_ ;
  assign \new_Sorter100|1645_  = \new_Sorter100|1544_  | \new_Sorter100|1545_ ;
  assign \new_Sorter100|1646_  = \new_Sorter100|1546_  & \new_Sorter100|1547_ ;
  assign \new_Sorter100|1647_  = \new_Sorter100|1546_  | \new_Sorter100|1547_ ;
  assign \new_Sorter100|1648_  = \new_Sorter100|1548_  & \new_Sorter100|1549_ ;
  assign \new_Sorter100|1649_  = \new_Sorter100|1548_  | \new_Sorter100|1549_ ;
  assign \new_Sorter100|1650_  = \new_Sorter100|1550_  & \new_Sorter100|1551_ ;
  assign \new_Sorter100|1651_  = \new_Sorter100|1550_  | \new_Sorter100|1551_ ;
  assign \new_Sorter100|1652_  = \new_Sorter100|1552_  & \new_Sorter100|1553_ ;
  assign \new_Sorter100|1653_  = \new_Sorter100|1552_  | \new_Sorter100|1553_ ;
  assign \new_Sorter100|1654_  = \new_Sorter100|1554_  & \new_Sorter100|1555_ ;
  assign \new_Sorter100|1655_  = \new_Sorter100|1554_  | \new_Sorter100|1555_ ;
  assign \new_Sorter100|1656_  = \new_Sorter100|1556_  & \new_Sorter100|1557_ ;
  assign \new_Sorter100|1657_  = \new_Sorter100|1556_  | \new_Sorter100|1557_ ;
  assign \new_Sorter100|1658_  = \new_Sorter100|1558_  & \new_Sorter100|1559_ ;
  assign \new_Sorter100|1659_  = \new_Sorter100|1558_  | \new_Sorter100|1559_ ;
  assign \new_Sorter100|1660_  = \new_Sorter100|1560_  & \new_Sorter100|1561_ ;
  assign \new_Sorter100|1661_  = \new_Sorter100|1560_  | \new_Sorter100|1561_ ;
  assign \new_Sorter100|1662_  = \new_Sorter100|1562_  & \new_Sorter100|1563_ ;
  assign \new_Sorter100|1663_  = \new_Sorter100|1562_  | \new_Sorter100|1563_ ;
  assign \new_Sorter100|1664_  = \new_Sorter100|1564_  & \new_Sorter100|1565_ ;
  assign \new_Sorter100|1665_  = \new_Sorter100|1564_  | \new_Sorter100|1565_ ;
  assign \new_Sorter100|1666_  = \new_Sorter100|1566_  & \new_Sorter100|1567_ ;
  assign \new_Sorter100|1667_  = \new_Sorter100|1566_  | \new_Sorter100|1567_ ;
  assign \new_Sorter100|1668_  = \new_Sorter100|1568_  & \new_Sorter100|1569_ ;
  assign \new_Sorter100|1669_  = \new_Sorter100|1568_  | \new_Sorter100|1569_ ;
  assign \new_Sorter100|1670_  = \new_Sorter100|1570_  & \new_Sorter100|1571_ ;
  assign \new_Sorter100|1671_  = \new_Sorter100|1570_  | \new_Sorter100|1571_ ;
  assign \new_Sorter100|1672_  = \new_Sorter100|1572_  & \new_Sorter100|1573_ ;
  assign \new_Sorter100|1673_  = \new_Sorter100|1572_  | \new_Sorter100|1573_ ;
  assign \new_Sorter100|1674_  = \new_Sorter100|1574_  & \new_Sorter100|1575_ ;
  assign \new_Sorter100|1675_  = \new_Sorter100|1574_  | \new_Sorter100|1575_ ;
  assign \new_Sorter100|1676_  = \new_Sorter100|1576_  & \new_Sorter100|1577_ ;
  assign \new_Sorter100|1677_  = \new_Sorter100|1576_  | \new_Sorter100|1577_ ;
  assign \new_Sorter100|1678_  = \new_Sorter100|1578_  & \new_Sorter100|1579_ ;
  assign \new_Sorter100|1679_  = \new_Sorter100|1578_  | \new_Sorter100|1579_ ;
  assign \new_Sorter100|1680_  = \new_Sorter100|1580_  & \new_Sorter100|1581_ ;
  assign \new_Sorter100|1681_  = \new_Sorter100|1580_  | \new_Sorter100|1581_ ;
  assign \new_Sorter100|1682_  = \new_Sorter100|1582_  & \new_Sorter100|1583_ ;
  assign \new_Sorter100|1683_  = \new_Sorter100|1582_  | \new_Sorter100|1583_ ;
  assign \new_Sorter100|1684_  = \new_Sorter100|1584_  & \new_Sorter100|1585_ ;
  assign \new_Sorter100|1685_  = \new_Sorter100|1584_  | \new_Sorter100|1585_ ;
  assign \new_Sorter100|1686_  = \new_Sorter100|1586_  & \new_Sorter100|1587_ ;
  assign \new_Sorter100|1687_  = \new_Sorter100|1586_  | \new_Sorter100|1587_ ;
  assign \new_Sorter100|1688_  = \new_Sorter100|1588_  & \new_Sorter100|1589_ ;
  assign \new_Sorter100|1689_  = \new_Sorter100|1588_  | \new_Sorter100|1589_ ;
  assign \new_Sorter100|1690_  = \new_Sorter100|1590_  & \new_Sorter100|1591_ ;
  assign \new_Sorter100|1691_  = \new_Sorter100|1590_  | \new_Sorter100|1591_ ;
  assign \new_Sorter100|1692_  = \new_Sorter100|1592_  & \new_Sorter100|1593_ ;
  assign \new_Sorter100|1693_  = \new_Sorter100|1592_  | \new_Sorter100|1593_ ;
  assign \new_Sorter100|1694_  = \new_Sorter100|1594_  & \new_Sorter100|1595_ ;
  assign \new_Sorter100|1695_  = \new_Sorter100|1594_  | \new_Sorter100|1595_ ;
  assign \new_Sorter100|1696_  = \new_Sorter100|1596_  & \new_Sorter100|1597_ ;
  assign \new_Sorter100|1697_  = \new_Sorter100|1596_  | \new_Sorter100|1597_ ;
  assign \new_Sorter100|1698_  = \new_Sorter100|1598_  & \new_Sorter100|1599_ ;
  assign \new_Sorter100|1699_  = \new_Sorter100|1598_  | \new_Sorter100|1599_ ;
  assign \new_Sorter100|1700_  = \new_Sorter100|1600_ ;
  assign \new_Sorter100|1799_  = \new_Sorter100|1699_ ;
  assign \new_Sorter100|1701_  = \new_Sorter100|1601_  & \new_Sorter100|1602_ ;
  assign \new_Sorter100|1702_  = \new_Sorter100|1601_  | \new_Sorter100|1602_ ;
  assign \new_Sorter100|1703_  = \new_Sorter100|1603_  & \new_Sorter100|1604_ ;
  assign \new_Sorter100|1704_  = \new_Sorter100|1603_  | \new_Sorter100|1604_ ;
  assign \new_Sorter100|1705_  = \new_Sorter100|1605_  & \new_Sorter100|1606_ ;
  assign \new_Sorter100|1706_  = \new_Sorter100|1605_  | \new_Sorter100|1606_ ;
  assign \new_Sorter100|1707_  = \new_Sorter100|1607_  & \new_Sorter100|1608_ ;
  assign \new_Sorter100|1708_  = \new_Sorter100|1607_  | \new_Sorter100|1608_ ;
  assign \new_Sorter100|1709_  = \new_Sorter100|1609_  & \new_Sorter100|1610_ ;
  assign \new_Sorter100|1710_  = \new_Sorter100|1609_  | \new_Sorter100|1610_ ;
  assign \new_Sorter100|1711_  = \new_Sorter100|1611_  & \new_Sorter100|1612_ ;
  assign \new_Sorter100|1712_  = \new_Sorter100|1611_  | \new_Sorter100|1612_ ;
  assign \new_Sorter100|1713_  = \new_Sorter100|1613_  & \new_Sorter100|1614_ ;
  assign \new_Sorter100|1714_  = \new_Sorter100|1613_  | \new_Sorter100|1614_ ;
  assign \new_Sorter100|1715_  = \new_Sorter100|1615_  & \new_Sorter100|1616_ ;
  assign \new_Sorter100|1716_  = \new_Sorter100|1615_  | \new_Sorter100|1616_ ;
  assign \new_Sorter100|1717_  = \new_Sorter100|1617_  & \new_Sorter100|1618_ ;
  assign \new_Sorter100|1718_  = \new_Sorter100|1617_  | \new_Sorter100|1618_ ;
  assign \new_Sorter100|1719_  = \new_Sorter100|1619_  & \new_Sorter100|1620_ ;
  assign \new_Sorter100|1720_  = \new_Sorter100|1619_  | \new_Sorter100|1620_ ;
  assign \new_Sorter100|1721_  = \new_Sorter100|1621_  & \new_Sorter100|1622_ ;
  assign \new_Sorter100|1722_  = \new_Sorter100|1621_  | \new_Sorter100|1622_ ;
  assign \new_Sorter100|1723_  = \new_Sorter100|1623_  & \new_Sorter100|1624_ ;
  assign \new_Sorter100|1724_  = \new_Sorter100|1623_  | \new_Sorter100|1624_ ;
  assign \new_Sorter100|1725_  = \new_Sorter100|1625_  & \new_Sorter100|1626_ ;
  assign \new_Sorter100|1726_  = \new_Sorter100|1625_  | \new_Sorter100|1626_ ;
  assign \new_Sorter100|1727_  = \new_Sorter100|1627_  & \new_Sorter100|1628_ ;
  assign \new_Sorter100|1728_  = \new_Sorter100|1627_  | \new_Sorter100|1628_ ;
  assign \new_Sorter100|1729_  = \new_Sorter100|1629_  & \new_Sorter100|1630_ ;
  assign \new_Sorter100|1730_  = \new_Sorter100|1629_  | \new_Sorter100|1630_ ;
  assign \new_Sorter100|1731_  = \new_Sorter100|1631_  & \new_Sorter100|1632_ ;
  assign \new_Sorter100|1732_  = \new_Sorter100|1631_  | \new_Sorter100|1632_ ;
  assign \new_Sorter100|1733_  = \new_Sorter100|1633_  & \new_Sorter100|1634_ ;
  assign \new_Sorter100|1734_  = \new_Sorter100|1633_  | \new_Sorter100|1634_ ;
  assign \new_Sorter100|1735_  = \new_Sorter100|1635_  & \new_Sorter100|1636_ ;
  assign \new_Sorter100|1736_  = \new_Sorter100|1635_  | \new_Sorter100|1636_ ;
  assign \new_Sorter100|1737_  = \new_Sorter100|1637_  & \new_Sorter100|1638_ ;
  assign \new_Sorter100|1738_  = \new_Sorter100|1637_  | \new_Sorter100|1638_ ;
  assign \new_Sorter100|1739_  = \new_Sorter100|1639_  & \new_Sorter100|1640_ ;
  assign \new_Sorter100|1740_  = \new_Sorter100|1639_  | \new_Sorter100|1640_ ;
  assign \new_Sorter100|1741_  = \new_Sorter100|1641_  & \new_Sorter100|1642_ ;
  assign \new_Sorter100|1742_  = \new_Sorter100|1641_  | \new_Sorter100|1642_ ;
  assign \new_Sorter100|1743_  = \new_Sorter100|1643_  & \new_Sorter100|1644_ ;
  assign \new_Sorter100|1744_  = \new_Sorter100|1643_  | \new_Sorter100|1644_ ;
  assign \new_Sorter100|1745_  = \new_Sorter100|1645_  & \new_Sorter100|1646_ ;
  assign \new_Sorter100|1746_  = \new_Sorter100|1645_  | \new_Sorter100|1646_ ;
  assign \new_Sorter100|1747_  = \new_Sorter100|1647_  & \new_Sorter100|1648_ ;
  assign \new_Sorter100|1748_  = \new_Sorter100|1647_  | \new_Sorter100|1648_ ;
  assign \new_Sorter100|1749_  = \new_Sorter100|1649_  & \new_Sorter100|1650_ ;
  assign \new_Sorter100|1750_  = \new_Sorter100|1649_  | \new_Sorter100|1650_ ;
  assign \new_Sorter100|1751_  = \new_Sorter100|1651_  & \new_Sorter100|1652_ ;
  assign \new_Sorter100|1752_  = \new_Sorter100|1651_  | \new_Sorter100|1652_ ;
  assign \new_Sorter100|1753_  = \new_Sorter100|1653_  & \new_Sorter100|1654_ ;
  assign \new_Sorter100|1754_  = \new_Sorter100|1653_  | \new_Sorter100|1654_ ;
  assign \new_Sorter100|1755_  = \new_Sorter100|1655_  & \new_Sorter100|1656_ ;
  assign \new_Sorter100|1756_  = \new_Sorter100|1655_  | \new_Sorter100|1656_ ;
  assign \new_Sorter100|1757_  = \new_Sorter100|1657_  & \new_Sorter100|1658_ ;
  assign \new_Sorter100|1758_  = \new_Sorter100|1657_  | \new_Sorter100|1658_ ;
  assign \new_Sorter100|1759_  = \new_Sorter100|1659_  & \new_Sorter100|1660_ ;
  assign \new_Sorter100|1760_  = \new_Sorter100|1659_  | \new_Sorter100|1660_ ;
  assign \new_Sorter100|1761_  = \new_Sorter100|1661_  & \new_Sorter100|1662_ ;
  assign \new_Sorter100|1762_  = \new_Sorter100|1661_  | \new_Sorter100|1662_ ;
  assign \new_Sorter100|1763_  = \new_Sorter100|1663_  & \new_Sorter100|1664_ ;
  assign \new_Sorter100|1764_  = \new_Sorter100|1663_  | \new_Sorter100|1664_ ;
  assign \new_Sorter100|1765_  = \new_Sorter100|1665_  & \new_Sorter100|1666_ ;
  assign \new_Sorter100|1766_  = \new_Sorter100|1665_  | \new_Sorter100|1666_ ;
  assign \new_Sorter100|1767_  = \new_Sorter100|1667_  & \new_Sorter100|1668_ ;
  assign \new_Sorter100|1768_  = \new_Sorter100|1667_  | \new_Sorter100|1668_ ;
  assign \new_Sorter100|1769_  = \new_Sorter100|1669_  & \new_Sorter100|1670_ ;
  assign \new_Sorter100|1770_  = \new_Sorter100|1669_  | \new_Sorter100|1670_ ;
  assign \new_Sorter100|1771_  = \new_Sorter100|1671_  & \new_Sorter100|1672_ ;
  assign \new_Sorter100|1772_  = \new_Sorter100|1671_  | \new_Sorter100|1672_ ;
  assign \new_Sorter100|1773_  = \new_Sorter100|1673_  & \new_Sorter100|1674_ ;
  assign \new_Sorter100|1774_  = \new_Sorter100|1673_  | \new_Sorter100|1674_ ;
  assign \new_Sorter100|1775_  = \new_Sorter100|1675_  & \new_Sorter100|1676_ ;
  assign \new_Sorter100|1776_  = \new_Sorter100|1675_  | \new_Sorter100|1676_ ;
  assign \new_Sorter100|1777_  = \new_Sorter100|1677_  & \new_Sorter100|1678_ ;
  assign \new_Sorter100|1778_  = \new_Sorter100|1677_  | \new_Sorter100|1678_ ;
  assign \new_Sorter100|1779_  = \new_Sorter100|1679_  & \new_Sorter100|1680_ ;
  assign \new_Sorter100|1780_  = \new_Sorter100|1679_  | \new_Sorter100|1680_ ;
  assign \new_Sorter100|1781_  = \new_Sorter100|1681_  & \new_Sorter100|1682_ ;
  assign \new_Sorter100|1782_  = \new_Sorter100|1681_  | \new_Sorter100|1682_ ;
  assign \new_Sorter100|1783_  = \new_Sorter100|1683_  & \new_Sorter100|1684_ ;
  assign \new_Sorter100|1784_  = \new_Sorter100|1683_  | \new_Sorter100|1684_ ;
  assign \new_Sorter100|1785_  = \new_Sorter100|1685_  & \new_Sorter100|1686_ ;
  assign \new_Sorter100|1786_  = \new_Sorter100|1685_  | \new_Sorter100|1686_ ;
  assign \new_Sorter100|1787_  = \new_Sorter100|1687_  & \new_Sorter100|1688_ ;
  assign \new_Sorter100|1788_  = \new_Sorter100|1687_  | \new_Sorter100|1688_ ;
  assign \new_Sorter100|1789_  = \new_Sorter100|1689_  & \new_Sorter100|1690_ ;
  assign \new_Sorter100|1790_  = \new_Sorter100|1689_  | \new_Sorter100|1690_ ;
  assign \new_Sorter100|1791_  = \new_Sorter100|1691_  & \new_Sorter100|1692_ ;
  assign \new_Sorter100|1792_  = \new_Sorter100|1691_  | \new_Sorter100|1692_ ;
  assign \new_Sorter100|1793_  = \new_Sorter100|1693_  & \new_Sorter100|1694_ ;
  assign \new_Sorter100|1794_  = \new_Sorter100|1693_  | \new_Sorter100|1694_ ;
  assign \new_Sorter100|1795_  = \new_Sorter100|1695_  & \new_Sorter100|1696_ ;
  assign \new_Sorter100|1796_  = \new_Sorter100|1695_  | \new_Sorter100|1696_ ;
  assign \new_Sorter100|1797_  = \new_Sorter100|1697_  & \new_Sorter100|1698_ ;
  assign \new_Sorter100|1798_  = \new_Sorter100|1697_  | \new_Sorter100|1698_ ;
  assign \new_Sorter100|1800_  = \new_Sorter100|1700_  & \new_Sorter100|1701_ ;
  assign \new_Sorter100|1801_  = \new_Sorter100|1700_  | \new_Sorter100|1701_ ;
  assign \new_Sorter100|1802_  = \new_Sorter100|1702_  & \new_Sorter100|1703_ ;
  assign \new_Sorter100|1803_  = \new_Sorter100|1702_  | \new_Sorter100|1703_ ;
  assign \new_Sorter100|1804_  = \new_Sorter100|1704_  & \new_Sorter100|1705_ ;
  assign \new_Sorter100|1805_  = \new_Sorter100|1704_  | \new_Sorter100|1705_ ;
  assign \new_Sorter100|1806_  = \new_Sorter100|1706_  & \new_Sorter100|1707_ ;
  assign \new_Sorter100|1807_  = \new_Sorter100|1706_  | \new_Sorter100|1707_ ;
  assign \new_Sorter100|1808_  = \new_Sorter100|1708_  & \new_Sorter100|1709_ ;
  assign \new_Sorter100|1809_  = \new_Sorter100|1708_  | \new_Sorter100|1709_ ;
  assign \new_Sorter100|1810_  = \new_Sorter100|1710_  & \new_Sorter100|1711_ ;
  assign \new_Sorter100|1811_  = \new_Sorter100|1710_  | \new_Sorter100|1711_ ;
  assign \new_Sorter100|1812_  = \new_Sorter100|1712_  & \new_Sorter100|1713_ ;
  assign \new_Sorter100|1813_  = \new_Sorter100|1712_  | \new_Sorter100|1713_ ;
  assign \new_Sorter100|1814_  = \new_Sorter100|1714_  & \new_Sorter100|1715_ ;
  assign \new_Sorter100|1815_  = \new_Sorter100|1714_  | \new_Sorter100|1715_ ;
  assign \new_Sorter100|1816_  = \new_Sorter100|1716_  & \new_Sorter100|1717_ ;
  assign \new_Sorter100|1817_  = \new_Sorter100|1716_  | \new_Sorter100|1717_ ;
  assign \new_Sorter100|1818_  = \new_Sorter100|1718_  & \new_Sorter100|1719_ ;
  assign \new_Sorter100|1819_  = \new_Sorter100|1718_  | \new_Sorter100|1719_ ;
  assign \new_Sorter100|1820_  = \new_Sorter100|1720_  & \new_Sorter100|1721_ ;
  assign \new_Sorter100|1821_  = \new_Sorter100|1720_  | \new_Sorter100|1721_ ;
  assign \new_Sorter100|1822_  = \new_Sorter100|1722_  & \new_Sorter100|1723_ ;
  assign \new_Sorter100|1823_  = \new_Sorter100|1722_  | \new_Sorter100|1723_ ;
  assign \new_Sorter100|1824_  = \new_Sorter100|1724_  & \new_Sorter100|1725_ ;
  assign \new_Sorter100|1825_  = \new_Sorter100|1724_  | \new_Sorter100|1725_ ;
  assign \new_Sorter100|1826_  = \new_Sorter100|1726_  & \new_Sorter100|1727_ ;
  assign \new_Sorter100|1827_  = \new_Sorter100|1726_  | \new_Sorter100|1727_ ;
  assign \new_Sorter100|1828_  = \new_Sorter100|1728_  & \new_Sorter100|1729_ ;
  assign \new_Sorter100|1829_  = \new_Sorter100|1728_  | \new_Sorter100|1729_ ;
  assign \new_Sorter100|1830_  = \new_Sorter100|1730_  & \new_Sorter100|1731_ ;
  assign \new_Sorter100|1831_  = \new_Sorter100|1730_  | \new_Sorter100|1731_ ;
  assign \new_Sorter100|1832_  = \new_Sorter100|1732_  & \new_Sorter100|1733_ ;
  assign \new_Sorter100|1833_  = \new_Sorter100|1732_  | \new_Sorter100|1733_ ;
  assign \new_Sorter100|1834_  = \new_Sorter100|1734_  & \new_Sorter100|1735_ ;
  assign \new_Sorter100|1835_  = \new_Sorter100|1734_  | \new_Sorter100|1735_ ;
  assign \new_Sorter100|1836_  = \new_Sorter100|1736_  & \new_Sorter100|1737_ ;
  assign \new_Sorter100|1837_  = \new_Sorter100|1736_  | \new_Sorter100|1737_ ;
  assign \new_Sorter100|1838_  = \new_Sorter100|1738_  & \new_Sorter100|1739_ ;
  assign \new_Sorter100|1839_  = \new_Sorter100|1738_  | \new_Sorter100|1739_ ;
  assign \new_Sorter100|1840_  = \new_Sorter100|1740_  & \new_Sorter100|1741_ ;
  assign \new_Sorter100|1841_  = \new_Sorter100|1740_  | \new_Sorter100|1741_ ;
  assign \new_Sorter100|1842_  = \new_Sorter100|1742_  & \new_Sorter100|1743_ ;
  assign \new_Sorter100|1843_  = \new_Sorter100|1742_  | \new_Sorter100|1743_ ;
  assign \new_Sorter100|1844_  = \new_Sorter100|1744_  & \new_Sorter100|1745_ ;
  assign \new_Sorter100|1845_  = \new_Sorter100|1744_  | \new_Sorter100|1745_ ;
  assign \new_Sorter100|1846_  = \new_Sorter100|1746_  & \new_Sorter100|1747_ ;
  assign \new_Sorter100|1847_  = \new_Sorter100|1746_  | \new_Sorter100|1747_ ;
  assign \new_Sorter100|1848_  = \new_Sorter100|1748_  & \new_Sorter100|1749_ ;
  assign \new_Sorter100|1849_  = \new_Sorter100|1748_  | \new_Sorter100|1749_ ;
  assign \new_Sorter100|1850_  = \new_Sorter100|1750_  & \new_Sorter100|1751_ ;
  assign \new_Sorter100|1851_  = \new_Sorter100|1750_  | \new_Sorter100|1751_ ;
  assign \new_Sorter100|1852_  = \new_Sorter100|1752_  & \new_Sorter100|1753_ ;
  assign \new_Sorter100|1853_  = \new_Sorter100|1752_  | \new_Sorter100|1753_ ;
  assign \new_Sorter100|1854_  = \new_Sorter100|1754_  & \new_Sorter100|1755_ ;
  assign \new_Sorter100|1855_  = \new_Sorter100|1754_  | \new_Sorter100|1755_ ;
  assign \new_Sorter100|1856_  = \new_Sorter100|1756_  & \new_Sorter100|1757_ ;
  assign \new_Sorter100|1857_  = \new_Sorter100|1756_  | \new_Sorter100|1757_ ;
  assign \new_Sorter100|1858_  = \new_Sorter100|1758_  & \new_Sorter100|1759_ ;
  assign \new_Sorter100|1859_  = \new_Sorter100|1758_  | \new_Sorter100|1759_ ;
  assign \new_Sorter100|1860_  = \new_Sorter100|1760_  & \new_Sorter100|1761_ ;
  assign \new_Sorter100|1861_  = \new_Sorter100|1760_  | \new_Sorter100|1761_ ;
  assign \new_Sorter100|1862_  = \new_Sorter100|1762_  & \new_Sorter100|1763_ ;
  assign \new_Sorter100|1863_  = \new_Sorter100|1762_  | \new_Sorter100|1763_ ;
  assign \new_Sorter100|1864_  = \new_Sorter100|1764_  & \new_Sorter100|1765_ ;
  assign \new_Sorter100|1865_  = \new_Sorter100|1764_  | \new_Sorter100|1765_ ;
  assign \new_Sorter100|1866_  = \new_Sorter100|1766_  & \new_Sorter100|1767_ ;
  assign \new_Sorter100|1867_  = \new_Sorter100|1766_  | \new_Sorter100|1767_ ;
  assign \new_Sorter100|1868_  = \new_Sorter100|1768_  & \new_Sorter100|1769_ ;
  assign \new_Sorter100|1869_  = \new_Sorter100|1768_  | \new_Sorter100|1769_ ;
  assign \new_Sorter100|1870_  = \new_Sorter100|1770_  & \new_Sorter100|1771_ ;
  assign \new_Sorter100|1871_  = \new_Sorter100|1770_  | \new_Sorter100|1771_ ;
  assign \new_Sorter100|1872_  = \new_Sorter100|1772_  & \new_Sorter100|1773_ ;
  assign \new_Sorter100|1873_  = \new_Sorter100|1772_  | \new_Sorter100|1773_ ;
  assign \new_Sorter100|1874_  = \new_Sorter100|1774_  & \new_Sorter100|1775_ ;
  assign \new_Sorter100|1875_  = \new_Sorter100|1774_  | \new_Sorter100|1775_ ;
  assign \new_Sorter100|1876_  = \new_Sorter100|1776_  & \new_Sorter100|1777_ ;
  assign \new_Sorter100|1877_  = \new_Sorter100|1776_  | \new_Sorter100|1777_ ;
  assign \new_Sorter100|1878_  = \new_Sorter100|1778_  & \new_Sorter100|1779_ ;
  assign \new_Sorter100|1879_  = \new_Sorter100|1778_  | \new_Sorter100|1779_ ;
  assign \new_Sorter100|1880_  = \new_Sorter100|1780_  & \new_Sorter100|1781_ ;
  assign \new_Sorter100|1881_  = \new_Sorter100|1780_  | \new_Sorter100|1781_ ;
  assign \new_Sorter100|1882_  = \new_Sorter100|1782_  & \new_Sorter100|1783_ ;
  assign \new_Sorter100|1883_  = \new_Sorter100|1782_  | \new_Sorter100|1783_ ;
  assign \new_Sorter100|1884_  = \new_Sorter100|1784_  & \new_Sorter100|1785_ ;
  assign \new_Sorter100|1885_  = \new_Sorter100|1784_  | \new_Sorter100|1785_ ;
  assign \new_Sorter100|1886_  = \new_Sorter100|1786_  & \new_Sorter100|1787_ ;
  assign \new_Sorter100|1887_  = \new_Sorter100|1786_  | \new_Sorter100|1787_ ;
  assign \new_Sorter100|1888_  = \new_Sorter100|1788_  & \new_Sorter100|1789_ ;
  assign \new_Sorter100|1889_  = \new_Sorter100|1788_  | \new_Sorter100|1789_ ;
  assign \new_Sorter100|1890_  = \new_Sorter100|1790_  & \new_Sorter100|1791_ ;
  assign \new_Sorter100|1891_  = \new_Sorter100|1790_  | \new_Sorter100|1791_ ;
  assign \new_Sorter100|1892_  = \new_Sorter100|1792_  & \new_Sorter100|1793_ ;
  assign \new_Sorter100|1893_  = \new_Sorter100|1792_  | \new_Sorter100|1793_ ;
  assign \new_Sorter100|1894_  = \new_Sorter100|1794_  & \new_Sorter100|1795_ ;
  assign \new_Sorter100|1895_  = \new_Sorter100|1794_  | \new_Sorter100|1795_ ;
  assign \new_Sorter100|1896_  = \new_Sorter100|1796_  & \new_Sorter100|1797_ ;
  assign \new_Sorter100|1897_  = \new_Sorter100|1796_  | \new_Sorter100|1797_ ;
  assign \new_Sorter100|1898_  = \new_Sorter100|1798_  & \new_Sorter100|1799_ ;
  assign \new_Sorter100|1899_  = \new_Sorter100|1798_  | \new_Sorter100|1799_ ;
  assign \new_Sorter100|1900_  = \new_Sorter100|1800_ ;
  assign \new_Sorter100|1999_  = \new_Sorter100|1899_ ;
  assign \new_Sorter100|1901_  = \new_Sorter100|1801_  & \new_Sorter100|1802_ ;
  assign \new_Sorter100|1902_  = \new_Sorter100|1801_  | \new_Sorter100|1802_ ;
  assign \new_Sorter100|1903_  = \new_Sorter100|1803_  & \new_Sorter100|1804_ ;
  assign \new_Sorter100|1904_  = \new_Sorter100|1803_  | \new_Sorter100|1804_ ;
  assign \new_Sorter100|1905_  = \new_Sorter100|1805_  & \new_Sorter100|1806_ ;
  assign \new_Sorter100|1906_  = \new_Sorter100|1805_  | \new_Sorter100|1806_ ;
  assign \new_Sorter100|1907_  = \new_Sorter100|1807_  & \new_Sorter100|1808_ ;
  assign \new_Sorter100|1908_  = \new_Sorter100|1807_  | \new_Sorter100|1808_ ;
  assign \new_Sorter100|1909_  = \new_Sorter100|1809_  & \new_Sorter100|1810_ ;
  assign \new_Sorter100|1910_  = \new_Sorter100|1809_  | \new_Sorter100|1810_ ;
  assign \new_Sorter100|1911_  = \new_Sorter100|1811_  & \new_Sorter100|1812_ ;
  assign \new_Sorter100|1912_  = \new_Sorter100|1811_  | \new_Sorter100|1812_ ;
  assign \new_Sorter100|1913_  = \new_Sorter100|1813_  & \new_Sorter100|1814_ ;
  assign \new_Sorter100|1914_  = \new_Sorter100|1813_  | \new_Sorter100|1814_ ;
  assign \new_Sorter100|1915_  = \new_Sorter100|1815_  & \new_Sorter100|1816_ ;
  assign \new_Sorter100|1916_  = \new_Sorter100|1815_  | \new_Sorter100|1816_ ;
  assign \new_Sorter100|1917_  = \new_Sorter100|1817_  & \new_Sorter100|1818_ ;
  assign \new_Sorter100|1918_  = \new_Sorter100|1817_  | \new_Sorter100|1818_ ;
  assign \new_Sorter100|1919_  = \new_Sorter100|1819_  & \new_Sorter100|1820_ ;
  assign \new_Sorter100|1920_  = \new_Sorter100|1819_  | \new_Sorter100|1820_ ;
  assign \new_Sorter100|1921_  = \new_Sorter100|1821_  & \new_Sorter100|1822_ ;
  assign \new_Sorter100|1922_  = \new_Sorter100|1821_  | \new_Sorter100|1822_ ;
  assign \new_Sorter100|1923_  = \new_Sorter100|1823_  & \new_Sorter100|1824_ ;
  assign \new_Sorter100|1924_  = \new_Sorter100|1823_  | \new_Sorter100|1824_ ;
  assign \new_Sorter100|1925_  = \new_Sorter100|1825_  & \new_Sorter100|1826_ ;
  assign \new_Sorter100|1926_  = \new_Sorter100|1825_  | \new_Sorter100|1826_ ;
  assign \new_Sorter100|1927_  = \new_Sorter100|1827_  & \new_Sorter100|1828_ ;
  assign \new_Sorter100|1928_  = \new_Sorter100|1827_  | \new_Sorter100|1828_ ;
  assign \new_Sorter100|1929_  = \new_Sorter100|1829_  & \new_Sorter100|1830_ ;
  assign \new_Sorter100|1930_  = \new_Sorter100|1829_  | \new_Sorter100|1830_ ;
  assign \new_Sorter100|1931_  = \new_Sorter100|1831_  & \new_Sorter100|1832_ ;
  assign \new_Sorter100|1932_  = \new_Sorter100|1831_  | \new_Sorter100|1832_ ;
  assign \new_Sorter100|1933_  = \new_Sorter100|1833_  & \new_Sorter100|1834_ ;
  assign \new_Sorter100|1934_  = \new_Sorter100|1833_  | \new_Sorter100|1834_ ;
  assign \new_Sorter100|1935_  = \new_Sorter100|1835_  & \new_Sorter100|1836_ ;
  assign \new_Sorter100|1936_  = \new_Sorter100|1835_  | \new_Sorter100|1836_ ;
  assign \new_Sorter100|1937_  = \new_Sorter100|1837_  & \new_Sorter100|1838_ ;
  assign \new_Sorter100|1938_  = \new_Sorter100|1837_  | \new_Sorter100|1838_ ;
  assign \new_Sorter100|1939_  = \new_Sorter100|1839_  & \new_Sorter100|1840_ ;
  assign \new_Sorter100|1940_  = \new_Sorter100|1839_  | \new_Sorter100|1840_ ;
  assign \new_Sorter100|1941_  = \new_Sorter100|1841_  & \new_Sorter100|1842_ ;
  assign \new_Sorter100|1942_  = \new_Sorter100|1841_  | \new_Sorter100|1842_ ;
  assign \new_Sorter100|1943_  = \new_Sorter100|1843_  & \new_Sorter100|1844_ ;
  assign \new_Sorter100|1944_  = \new_Sorter100|1843_  | \new_Sorter100|1844_ ;
  assign \new_Sorter100|1945_  = \new_Sorter100|1845_  & \new_Sorter100|1846_ ;
  assign \new_Sorter100|1946_  = \new_Sorter100|1845_  | \new_Sorter100|1846_ ;
  assign \new_Sorter100|1947_  = \new_Sorter100|1847_  & \new_Sorter100|1848_ ;
  assign \new_Sorter100|1948_  = \new_Sorter100|1847_  | \new_Sorter100|1848_ ;
  assign \new_Sorter100|1949_  = \new_Sorter100|1849_  & \new_Sorter100|1850_ ;
  assign \new_Sorter100|1950_  = \new_Sorter100|1849_  | \new_Sorter100|1850_ ;
  assign \new_Sorter100|1951_  = \new_Sorter100|1851_  & \new_Sorter100|1852_ ;
  assign \new_Sorter100|1952_  = \new_Sorter100|1851_  | \new_Sorter100|1852_ ;
  assign \new_Sorter100|1953_  = \new_Sorter100|1853_  & \new_Sorter100|1854_ ;
  assign \new_Sorter100|1954_  = \new_Sorter100|1853_  | \new_Sorter100|1854_ ;
  assign \new_Sorter100|1955_  = \new_Sorter100|1855_  & \new_Sorter100|1856_ ;
  assign \new_Sorter100|1956_  = \new_Sorter100|1855_  | \new_Sorter100|1856_ ;
  assign \new_Sorter100|1957_  = \new_Sorter100|1857_  & \new_Sorter100|1858_ ;
  assign \new_Sorter100|1958_  = \new_Sorter100|1857_  | \new_Sorter100|1858_ ;
  assign \new_Sorter100|1959_  = \new_Sorter100|1859_  & \new_Sorter100|1860_ ;
  assign \new_Sorter100|1960_  = \new_Sorter100|1859_  | \new_Sorter100|1860_ ;
  assign \new_Sorter100|1961_  = \new_Sorter100|1861_  & \new_Sorter100|1862_ ;
  assign \new_Sorter100|1962_  = \new_Sorter100|1861_  | \new_Sorter100|1862_ ;
  assign \new_Sorter100|1963_  = \new_Sorter100|1863_  & \new_Sorter100|1864_ ;
  assign \new_Sorter100|1964_  = \new_Sorter100|1863_  | \new_Sorter100|1864_ ;
  assign \new_Sorter100|1965_  = \new_Sorter100|1865_  & \new_Sorter100|1866_ ;
  assign \new_Sorter100|1966_  = \new_Sorter100|1865_  | \new_Sorter100|1866_ ;
  assign \new_Sorter100|1967_  = \new_Sorter100|1867_  & \new_Sorter100|1868_ ;
  assign \new_Sorter100|1968_  = \new_Sorter100|1867_  | \new_Sorter100|1868_ ;
  assign \new_Sorter100|1969_  = \new_Sorter100|1869_  & \new_Sorter100|1870_ ;
  assign \new_Sorter100|1970_  = \new_Sorter100|1869_  | \new_Sorter100|1870_ ;
  assign \new_Sorter100|1971_  = \new_Sorter100|1871_  & \new_Sorter100|1872_ ;
  assign \new_Sorter100|1972_  = \new_Sorter100|1871_  | \new_Sorter100|1872_ ;
  assign \new_Sorter100|1973_  = \new_Sorter100|1873_  & \new_Sorter100|1874_ ;
  assign \new_Sorter100|1974_  = \new_Sorter100|1873_  | \new_Sorter100|1874_ ;
  assign \new_Sorter100|1975_  = \new_Sorter100|1875_  & \new_Sorter100|1876_ ;
  assign \new_Sorter100|1976_  = \new_Sorter100|1875_  | \new_Sorter100|1876_ ;
  assign \new_Sorter100|1977_  = \new_Sorter100|1877_  & \new_Sorter100|1878_ ;
  assign \new_Sorter100|1978_  = \new_Sorter100|1877_  | \new_Sorter100|1878_ ;
  assign \new_Sorter100|1979_  = \new_Sorter100|1879_  & \new_Sorter100|1880_ ;
  assign \new_Sorter100|1980_  = \new_Sorter100|1879_  | \new_Sorter100|1880_ ;
  assign \new_Sorter100|1981_  = \new_Sorter100|1881_  & \new_Sorter100|1882_ ;
  assign \new_Sorter100|1982_  = \new_Sorter100|1881_  | \new_Sorter100|1882_ ;
  assign \new_Sorter100|1983_  = \new_Sorter100|1883_  & \new_Sorter100|1884_ ;
  assign \new_Sorter100|1984_  = \new_Sorter100|1883_  | \new_Sorter100|1884_ ;
  assign \new_Sorter100|1985_  = \new_Sorter100|1885_  & \new_Sorter100|1886_ ;
  assign \new_Sorter100|1986_  = \new_Sorter100|1885_  | \new_Sorter100|1886_ ;
  assign \new_Sorter100|1987_  = \new_Sorter100|1887_  & \new_Sorter100|1888_ ;
  assign \new_Sorter100|1988_  = \new_Sorter100|1887_  | \new_Sorter100|1888_ ;
  assign \new_Sorter100|1989_  = \new_Sorter100|1889_  & \new_Sorter100|1890_ ;
  assign \new_Sorter100|1990_  = \new_Sorter100|1889_  | \new_Sorter100|1890_ ;
  assign \new_Sorter100|1991_  = \new_Sorter100|1891_  & \new_Sorter100|1892_ ;
  assign \new_Sorter100|1992_  = \new_Sorter100|1891_  | \new_Sorter100|1892_ ;
  assign \new_Sorter100|1993_  = \new_Sorter100|1893_  & \new_Sorter100|1894_ ;
  assign \new_Sorter100|1994_  = \new_Sorter100|1893_  | \new_Sorter100|1894_ ;
  assign \new_Sorter100|1995_  = \new_Sorter100|1895_  & \new_Sorter100|1896_ ;
  assign \new_Sorter100|1996_  = \new_Sorter100|1895_  | \new_Sorter100|1896_ ;
  assign \new_Sorter100|1997_  = \new_Sorter100|1897_  & \new_Sorter100|1898_ ;
  assign \new_Sorter100|1998_  = \new_Sorter100|1897_  | \new_Sorter100|1898_ ;
  assign \new_Sorter100|2000_  = \new_Sorter100|1900_  & \new_Sorter100|1901_ ;
  assign \new_Sorter100|2001_  = \new_Sorter100|1900_  | \new_Sorter100|1901_ ;
  assign \new_Sorter100|2002_  = \new_Sorter100|1902_  & \new_Sorter100|1903_ ;
  assign \new_Sorter100|2003_  = \new_Sorter100|1902_  | \new_Sorter100|1903_ ;
  assign \new_Sorter100|2004_  = \new_Sorter100|1904_  & \new_Sorter100|1905_ ;
  assign \new_Sorter100|2005_  = \new_Sorter100|1904_  | \new_Sorter100|1905_ ;
  assign \new_Sorter100|2006_  = \new_Sorter100|1906_  & \new_Sorter100|1907_ ;
  assign \new_Sorter100|2007_  = \new_Sorter100|1906_  | \new_Sorter100|1907_ ;
  assign \new_Sorter100|2008_  = \new_Sorter100|1908_  & \new_Sorter100|1909_ ;
  assign \new_Sorter100|2009_  = \new_Sorter100|1908_  | \new_Sorter100|1909_ ;
  assign \new_Sorter100|2010_  = \new_Sorter100|1910_  & \new_Sorter100|1911_ ;
  assign \new_Sorter100|2011_  = \new_Sorter100|1910_  | \new_Sorter100|1911_ ;
  assign \new_Sorter100|2012_  = \new_Sorter100|1912_  & \new_Sorter100|1913_ ;
  assign \new_Sorter100|2013_  = \new_Sorter100|1912_  | \new_Sorter100|1913_ ;
  assign \new_Sorter100|2014_  = \new_Sorter100|1914_  & \new_Sorter100|1915_ ;
  assign \new_Sorter100|2015_  = \new_Sorter100|1914_  | \new_Sorter100|1915_ ;
  assign \new_Sorter100|2016_  = \new_Sorter100|1916_  & \new_Sorter100|1917_ ;
  assign \new_Sorter100|2017_  = \new_Sorter100|1916_  | \new_Sorter100|1917_ ;
  assign \new_Sorter100|2018_  = \new_Sorter100|1918_  & \new_Sorter100|1919_ ;
  assign \new_Sorter100|2019_  = \new_Sorter100|1918_  | \new_Sorter100|1919_ ;
  assign \new_Sorter100|2020_  = \new_Sorter100|1920_  & \new_Sorter100|1921_ ;
  assign \new_Sorter100|2021_  = \new_Sorter100|1920_  | \new_Sorter100|1921_ ;
  assign \new_Sorter100|2022_  = \new_Sorter100|1922_  & \new_Sorter100|1923_ ;
  assign \new_Sorter100|2023_  = \new_Sorter100|1922_  | \new_Sorter100|1923_ ;
  assign \new_Sorter100|2024_  = \new_Sorter100|1924_  & \new_Sorter100|1925_ ;
  assign \new_Sorter100|2025_  = \new_Sorter100|1924_  | \new_Sorter100|1925_ ;
  assign \new_Sorter100|2026_  = \new_Sorter100|1926_  & \new_Sorter100|1927_ ;
  assign \new_Sorter100|2027_  = \new_Sorter100|1926_  | \new_Sorter100|1927_ ;
  assign \new_Sorter100|2028_  = \new_Sorter100|1928_  & \new_Sorter100|1929_ ;
  assign \new_Sorter100|2029_  = \new_Sorter100|1928_  | \new_Sorter100|1929_ ;
  assign \new_Sorter100|2030_  = \new_Sorter100|1930_  & \new_Sorter100|1931_ ;
  assign \new_Sorter100|2031_  = \new_Sorter100|1930_  | \new_Sorter100|1931_ ;
  assign \new_Sorter100|2032_  = \new_Sorter100|1932_  & \new_Sorter100|1933_ ;
  assign \new_Sorter100|2033_  = \new_Sorter100|1932_  | \new_Sorter100|1933_ ;
  assign \new_Sorter100|2034_  = \new_Sorter100|1934_  & \new_Sorter100|1935_ ;
  assign \new_Sorter100|2035_  = \new_Sorter100|1934_  | \new_Sorter100|1935_ ;
  assign \new_Sorter100|2036_  = \new_Sorter100|1936_  & \new_Sorter100|1937_ ;
  assign \new_Sorter100|2037_  = \new_Sorter100|1936_  | \new_Sorter100|1937_ ;
  assign \new_Sorter100|2038_  = \new_Sorter100|1938_  & \new_Sorter100|1939_ ;
  assign \new_Sorter100|2039_  = \new_Sorter100|1938_  | \new_Sorter100|1939_ ;
  assign \new_Sorter100|2040_  = \new_Sorter100|1940_  & \new_Sorter100|1941_ ;
  assign \new_Sorter100|2041_  = \new_Sorter100|1940_  | \new_Sorter100|1941_ ;
  assign \new_Sorter100|2042_  = \new_Sorter100|1942_  & \new_Sorter100|1943_ ;
  assign \new_Sorter100|2043_  = \new_Sorter100|1942_  | \new_Sorter100|1943_ ;
  assign \new_Sorter100|2044_  = \new_Sorter100|1944_  & \new_Sorter100|1945_ ;
  assign \new_Sorter100|2045_  = \new_Sorter100|1944_  | \new_Sorter100|1945_ ;
  assign \new_Sorter100|2046_  = \new_Sorter100|1946_  & \new_Sorter100|1947_ ;
  assign \new_Sorter100|2047_  = \new_Sorter100|1946_  | \new_Sorter100|1947_ ;
  assign \new_Sorter100|2048_  = \new_Sorter100|1948_  & \new_Sorter100|1949_ ;
  assign \new_Sorter100|2049_  = \new_Sorter100|1948_  | \new_Sorter100|1949_ ;
  assign \new_Sorter100|2050_  = \new_Sorter100|1950_  & \new_Sorter100|1951_ ;
  assign \new_Sorter100|2051_  = \new_Sorter100|1950_  | \new_Sorter100|1951_ ;
  assign \new_Sorter100|2052_  = \new_Sorter100|1952_  & \new_Sorter100|1953_ ;
  assign \new_Sorter100|2053_  = \new_Sorter100|1952_  | \new_Sorter100|1953_ ;
  assign \new_Sorter100|2054_  = \new_Sorter100|1954_  & \new_Sorter100|1955_ ;
  assign \new_Sorter100|2055_  = \new_Sorter100|1954_  | \new_Sorter100|1955_ ;
  assign \new_Sorter100|2056_  = \new_Sorter100|1956_  & \new_Sorter100|1957_ ;
  assign \new_Sorter100|2057_  = \new_Sorter100|1956_  | \new_Sorter100|1957_ ;
  assign \new_Sorter100|2058_  = \new_Sorter100|1958_  & \new_Sorter100|1959_ ;
  assign \new_Sorter100|2059_  = \new_Sorter100|1958_  | \new_Sorter100|1959_ ;
  assign \new_Sorter100|2060_  = \new_Sorter100|1960_  & \new_Sorter100|1961_ ;
  assign \new_Sorter100|2061_  = \new_Sorter100|1960_  | \new_Sorter100|1961_ ;
  assign \new_Sorter100|2062_  = \new_Sorter100|1962_  & \new_Sorter100|1963_ ;
  assign \new_Sorter100|2063_  = \new_Sorter100|1962_  | \new_Sorter100|1963_ ;
  assign \new_Sorter100|2064_  = \new_Sorter100|1964_  & \new_Sorter100|1965_ ;
  assign \new_Sorter100|2065_  = \new_Sorter100|1964_  | \new_Sorter100|1965_ ;
  assign \new_Sorter100|2066_  = \new_Sorter100|1966_  & \new_Sorter100|1967_ ;
  assign \new_Sorter100|2067_  = \new_Sorter100|1966_  | \new_Sorter100|1967_ ;
  assign \new_Sorter100|2068_  = \new_Sorter100|1968_  & \new_Sorter100|1969_ ;
  assign \new_Sorter100|2069_  = \new_Sorter100|1968_  | \new_Sorter100|1969_ ;
  assign \new_Sorter100|2070_  = \new_Sorter100|1970_  & \new_Sorter100|1971_ ;
  assign \new_Sorter100|2071_  = \new_Sorter100|1970_  | \new_Sorter100|1971_ ;
  assign \new_Sorter100|2072_  = \new_Sorter100|1972_  & \new_Sorter100|1973_ ;
  assign \new_Sorter100|2073_  = \new_Sorter100|1972_  | \new_Sorter100|1973_ ;
  assign \new_Sorter100|2074_  = \new_Sorter100|1974_  & \new_Sorter100|1975_ ;
  assign \new_Sorter100|2075_  = \new_Sorter100|1974_  | \new_Sorter100|1975_ ;
  assign \new_Sorter100|2076_  = \new_Sorter100|1976_  & \new_Sorter100|1977_ ;
  assign \new_Sorter100|2077_  = \new_Sorter100|1976_  | \new_Sorter100|1977_ ;
  assign \new_Sorter100|2078_  = \new_Sorter100|1978_  & \new_Sorter100|1979_ ;
  assign \new_Sorter100|2079_  = \new_Sorter100|1978_  | \new_Sorter100|1979_ ;
  assign \new_Sorter100|2080_  = \new_Sorter100|1980_  & \new_Sorter100|1981_ ;
  assign \new_Sorter100|2081_  = \new_Sorter100|1980_  | \new_Sorter100|1981_ ;
  assign \new_Sorter100|2082_  = \new_Sorter100|1982_  & \new_Sorter100|1983_ ;
  assign \new_Sorter100|2083_  = \new_Sorter100|1982_  | \new_Sorter100|1983_ ;
  assign \new_Sorter100|2084_  = \new_Sorter100|1984_  & \new_Sorter100|1985_ ;
  assign \new_Sorter100|2085_  = \new_Sorter100|1984_  | \new_Sorter100|1985_ ;
  assign \new_Sorter100|2086_  = \new_Sorter100|1986_  & \new_Sorter100|1987_ ;
  assign \new_Sorter100|2087_  = \new_Sorter100|1986_  | \new_Sorter100|1987_ ;
  assign \new_Sorter100|2088_  = \new_Sorter100|1988_  & \new_Sorter100|1989_ ;
  assign \new_Sorter100|2089_  = \new_Sorter100|1988_  | \new_Sorter100|1989_ ;
  assign \new_Sorter100|2090_  = \new_Sorter100|1990_  & \new_Sorter100|1991_ ;
  assign \new_Sorter100|2091_  = \new_Sorter100|1990_  | \new_Sorter100|1991_ ;
  assign \new_Sorter100|2092_  = \new_Sorter100|1992_  & \new_Sorter100|1993_ ;
  assign \new_Sorter100|2093_  = \new_Sorter100|1992_  | \new_Sorter100|1993_ ;
  assign \new_Sorter100|2094_  = \new_Sorter100|1994_  & \new_Sorter100|1995_ ;
  assign \new_Sorter100|2095_  = \new_Sorter100|1994_  | \new_Sorter100|1995_ ;
  assign \new_Sorter100|2096_  = \new_Sorter100|1996_  & \new_Sorter100|1997_ ;
  assign \new_Sorter100|2097_  = \new_Sorter100|1996_  | \new_Sorter100|1997_ ;
  assign \new_Sorter100|2098_  = \new_Sorter100|1998_  & \new_Sorter100|1999_ ;
  assign \new_Sorter100|2099_  = \new_Sorter100|1998_  | \new_Sorter100|1999_ ;
  assign \new_Sorter100|2100_  = \new_Sorter100|2000_ ;
  assign \new_Sorter100|2199_  = \new_Sorter100|2099_ ;
  assign \new_Sorter100|2101_  = \new_Sorter100|2001_  & \new_Sorter100|2002_ ;
  assign \new_Sorter100|2102_  = \new_Sorter100|2001_  | \new_Sorter100|2002_ ;
  assign \new_Sorter100|2103_  = \new_Sorter100|2003_  & \new_Sorter100|2004_ ;
  assign \new_Sorter100|2104_  = \new_Sorter100|2003_  | \new_Sorter100|2004_ ;
  assign \new_Sorter100|2105_  = \new_Sorter100|2005_  & \new_Sorter100|2006_ ;
  assign \new_Sorter100|2106_  = \new_Sorter100|2005_  | \new_Sorter100|2006_ ;
  assign \new_Sorter100|2107_  = \new_Sorter100|2007_  & \new_Sorter100|2008_ ;
  assign \new_Sorter100|2108_  = \new_Sorter100|2007_  | \new_Sorter100|2008_ ;
  assign \new_Sorter100|2109_  = \new_Sorter100|2009_  & \new_Sorter100|2010_ ;
  assign \new_Sorter100|2110_  = \new_Sorter100|2009_  | \new_Sorter100|2010_ ;
  assign \new_Sorter100|2111_  = \new_Sorter100|2011_  & \new_Sorter100|2012_ ;
  assign \new_Sorter100|2112_  = \new_Sorter100|2011_  | \new_Sorter100|2012_ ;
  assign \new_Sorter100|2113_  = \new_Sorter100|2013_  & \new_Sorter100|2014_ ;
  assign \new_Sorter100|2114_  = \new_Sorter100|2013_  | \new_Sorter100|2014_ ;
  assign \new_Sorter100|2115_  = \new_Sorter100|2015_  & \new_Sorter100|2016_ ;
  assign \new_Sorter100|2116_  = \new_Sorter100|2015_  | \new_Sorter100|2016_ ;
  assign \new_Sorter100|2117_  = \new_Sorter100|2017_  & \new_Sorter100|2018_ ;
  assign \new_Sorter100|2118_  = \new_Sorter100|2017_  | \new_Sorter100|2018_ ;
  assign \new_Sorter100|2119_  = \new_Sorter100|2019_  & \new_Sorter100|2020_ ;
  assign \new_Sorter100|2120_  = \new_Sorter100|2019_  | \new_Sorter100|2020_ ;
  assign \new_Sorter100|2121_  = \new_Sorter100|2021_  & \new_Sorter100|2022_ ;
  assign \new_Sorter100|2122_  = \new_Sorter100|2021_  | \new_Sorter100|2022_ ;
  assign \new_Sorter100|2123_  = \new_Sorter100|2023_  & \new_Sorter100|2024_ ;
  assign \new_Sorter100|2124_  = \new_Sorter100|2023_  | \new_Sorter100|2024_ ;
  assign \new_Sorter100|2125_  = \new_Sorter100|2025_  & \new_Sorter100|2026_ ;
  assign \new_Sorter100|2126_  = \new_Sorter100|2025_  | \new_Sorter100|2026_ ;
  assign \new_Sorter100|2127_  = \new_Sorter100|2027_  & \new_Sorter100|2028_ ;
  assign \new_Sorter100|2128_  = \new_Sorter100|2027_  | \new_Sorter100|2028_ ;
  assign \new_Sorter100|2129_  = \new_Sorter100|2029_  & \new_Sorter100|2030_ ;
  assign \new_Sorter100|2130_  = \new_Sorter100|2029_  | \new_Sorter100|2030_ ;
  assign \new_Sorter100|2131_  = \new_Sorter100|2031_  & \new_Sorter100|2032_ ;
  assign \new_Sorter100|2132_  = \new_Sorter100|2031_  | \new_Sorter100|2032_ ;
  assign \new_Sorter100|2133_  = \new_Sorter100|2033_  & \new_Sorter100|2034_ ;
  assign \new_Sorter100|2134_  = \new_Sorter100|2033_  | \new_Sorter100|2034_ ;
  assign \new_Sorter100|2135_  = \new_Sorter100|2035_  & \new_Sorter100|2036_ ;
  assign \new_Sorter100|2136_  = \new_Sorter100|2035_  | \new_Sorter100|2036_ ;
  assign \new_Sorter100|2137_  = \new_Sorter100|2037_  & \new_Sorter100|2038_ ;
  assign \new_Sorter100|2138_  = \new_Sorter100|2037_  | \new_Sorter100|2038_ ;
  assign \new_Sorter100|2139_  = \new_Sorter100|2039_  & \new_Sorter100|2040_ ;
  assign \new_Sorter100|2140_  = \new_Sorter100|2039_  | \new_Sorter100|2040_ ;
  assign \new_Sorter100|2141_  = \new_Sorter100|2041_  & \new_Sorter100|2042_ ;
  assign \new_Sorter100|2142_  = \new_Sorter100|2041_  | \new_Sorter100|2042_ ;
  assign \new_Sorter100|2143_  = \new_Sorter100|2043_  & \new_Sorter100|2044_ ;
  assign \new_Sorter100|2144_  = \new_Sorter100|2043_  | \new_Sorter100|2044_ ;
  assign \new_Sorter100|2145_  = \new_Sorter100|2045_  & \new_Sorter100|2046_ ;
  assign \new_Sorter100|2146_  = \new_Sorter100|2045_  | \new_Sorter100|2046_ ;
  assign \new_Sorter100|2147_  = \new_Sorter100|2047_  & \new_Sorter100|2048_ ;
  assign \new_Sorter100|2148_  = \new_Sorter100|2047_  | \new_Sorter100|2048_ ;
  assign \new_Sorter100|2149_  = \new_Sorter100|2049_  & \new_Sorter100|2050_ ;
  assign \new_Sorter100|2150_  = \new_Sorter100|2049_  | \new_Sorter100|2050_ ;
  assign \new_Sorter100|2151_  = \new_Sorter100|2051_  & \new_Sorter100|2052_ ;
  assign \new_Sorter100|2152_  = \new_Sorter100|2051_  | \new_Sorter100|2052_ ;
  assign \new_Sorter100|2153_  = \new_Sorter100|2053_  & \new_Sorter100|2054_ ;
  assign \new_Sorter100|2154_  = \new_Sorter100|2053_  | \new_Sorter100|2054_ ;
  assign \new_Sorter100|2155_  = \new_Sorter100|2055_  & \new_Sorter100|2056_ ;
  assign \new_Sorter100|2156_  = \new_Sorter100|2055_  | \new_Sorter100|2056_ ;
  assign \new_Sorter100|2157_  = \new_Sorter100|2057_  & \new_Sorter100|2058_ ;
  assign \new_Sorter100|2158_  = \new_Sorter100|2057_  | \new_Sorter100|2058_ ;
  assign \new_Sorter100|2159_  = \new_Sorter100|2059_  & \new_Sorter100|2060_ ;
  assign \new_Sorter100|2160_  = \new_Sorter100|2059_  | \new_Sorter100|2060_ ;
  assign \new_Sorter100|2161_  = \new_Sorter100|2061_  & \new_Sorter100|2062_ ;
  assign \new_Sorter100|2162_  = \new_Sorter100|2061_  | \new_Sorter100|2062_ ;
  assign \new_Sorter100|2163_  = \new_Sorter100|2063_  & \new_Sorter100|2064_ ;
  assign \new_Sorter100|2164_  = \new_Sorter100|2063_  | \new_Sorter100|2064_ ;
  assign \new_Sorter100|2165_  = \new_Sorter100|2065_  & \new_Sorter100|2066_ ;
  assign \new_Sorter100|2166_  = \new_Sorter100|2065_  | \new_Sorter100|2066_ ;
  assign \new_Sorter100|2167_  = \new_Sorter100|2067_  & \new_Sorter100|2068_ ;
  assign \new_Sorter100|2168_  = \new_Sorter100|2067_  | \new_Sorter100|2068_ ;
  assign \new_Sorter100|2169_  = \new_Sorter100|2069_  & \new_Sorter100|2070_ ;
  assign \new_Sorter100|2170_  = \new_Sorter100|2069_  | \new_Sorter100|2070_ ;
  assign \new_Sorter100|2171_  = \new_Sorter100|2071_  & \new_Sorter100|2072_ ;
  assign \new_Sorter100|2172_  = \new_Sorter100|2071_  | \new_Sorter100|2072_ ;
  assign \new_Sorter100|2173_  = \new_Sorter100|2073_  & \new_Sorter100|2074_ ;
  assign \new_Sorter100|2174_  = \new_Sorter100|2073_  | \new_Sorter100|2074_ ;
  assign \new_Sorter100|2175_  = \new_Sorter100|2075_  & \new_Sorter100|2076_ ;
  assign \new_Sorter100|2176_  = \new_Sorter100|2075_  | \new_Sorter100|2076_ ;
  assign \new_Sorter100|2177_  = \new_Sorter100|2077_  & \new_Sorter100|2078_ ;
  assign \new_Sorter100|2178_  = \new_Sorter100|2077_  | \new_Sorter100|2078_ ;
  assign \new_Sorter100|2179_  = \new_Sorter100|2079_  & \new_Sorter100|2080_ ;
  assign \new_Sorter100|2180_  = \new_Sorter100|2079_  | \new_Sorter100|2080_ ;
  assign \new_Sorter100|2181_  = \new_Sorter100|2081_  & \new_Sorter100|2082_ ;
  assign \new_Sorter100|2182_  = \new_Sorter100|2081_  | \new_Sorter100|2082_ ;
  assign \new_Sorter100|2183_  = \new_Sorter100|2083_  & \new_Sorter100|2084_ ;
  assign \new_Sorter100|2184_  = \new_Sorter100|2083_  | \new_Sorter100|2084_ ;
  assign \new_Sorter100|2185_  = \new_Sorter100|2085_  & \new_Sorter100|2086_ ;
  assign \new_Sorter100|2186_  = \new_Sorter100|2085_  | \new_Sorter100|2086_ ;
  assign \new_Sorter100|2187_  = \new_Sorter100|2087_  & \new_Sorter100|2088_ ;
  assign \new_Sorter100|2188_  = \new_Sorter100|2087_  | \new_Sorter100|2088_ ;
  assign \new_Sorter100|2189_  = \new_Sorter100|2089_  & \new_Sorter100|2090_ ;
  assign \new_Sorter100|2190_  = \new_Sorter100|2089_  | \new_Sorter100|2090_ ;
  assign \new_Sorter100|2191_  = \new_Sorter100|2091_  & \new_Sorter100|2092_ ;
  assign \new_Sorter100|2192_  = \new_Sorter100|2091_  | \new_Sorter100|2092_ ;
  assign \new_Sorter100|2193_  = \new_Sorter100|2093_  & \new_Sorter100|2094_ ;
  assign \new_Sorter100|2194_  = \new_Sorter100|2093_  | \new_Sorter100|2094_ ;
  assign \new_Sorter100|2195_  = \new_Sorter100|2095_  & \new_Sorter100|2096_ ;
  assign \new_Sorter100|2196_  = \new_Sorter100|2095_  | \new_Sorter100|2096_ ;
  assign \new_Sorter100|2197_  = \new_Sorter100|2097_  & \new_Sorter100|2098_ ;
  assign \new_Sorter100|2198_  = \new_Sorter100|2097_  | \new_Sorter100|2098_ ;
  assign \new_Sorter100|2200_  = \new_Sorter100|2100_  & \new_Sorter100|2101_ ;
  assign \new_Sorter100|2201_  = \new_Sorter100|2100_  | \new_Sorter100|2101_ ;
  assign \new_Sorter100|2202_  = \new_Sorter100|2102_  & \new_Sorter100|2103_ ;
  assign \new_Sorter100|2203_  = \new_Sorter100|2102_  | \new_Sorter100|2103_ ;
  assign \new_Sorter100|2204_  = \new_Sorter100|2104_  & \new_Sorter100|2105_ ;
  assign \new_Sorter100|2205_  = \new_Sorter100|2104_  | \new_Sorter100|2105_ ;
  assign \new_Sorter100|2206_  = \new_Sorter100|2106_  & \new_Sorter100|2107_ ;
  assign \new_Sorter100|2207_  = \new_Sorter100|2106_  | \new_Sorter100|2107_ ;
  assign \new_Sorter100|2208_  = \new_Sorter100|2108_  & \new_Sorter100|2109_ ;
  assign \new_Sorter100|2209_  = \new_Sorter100|2108_  | \new_Sorter100|2109_ ;
  assign \new_Sorter100|2210_  = \new_Sorter100|2110_  & \new_Sorter100|2111_ ;
  assign \new_Sorter100|2211_  = \new_Sorter100|2110_  | \new_Sorter100|2111_ ;
  assign \new_Sorter100|2212_  = \new_Sorter100|2112_  & \new_Sorter100|2113_ ;
  assign \new_Sorter100|2213_  = \new_Sorter100|2112_  | \new_Sorter100|2113_ ;
  assign \new_Sorter100|2214_  = \new_Sorter100|2114_  & \new_Sorter100|2115_ ;
  assign \new_Sorter100|2215_  = \new_Sorter100|2114_  | \new_Sorter100|2115_ ;
  assign \new_Sorter100|2216_  = \new_Sorter100|2116_  & \new_Sorter100|2117_ ;
  assign \new_Sorter100|2217_  = \new_Sorter100|2116_  | \new_Sorter100|2117_ ;
  assign \new_Sorter100|2218_  = \new_Sorter100|2118_  & \new_Sorter100|2119_ ;
  assign \new_Sorter100|2219_  = \new_Sorter100|2118_  | \new_Sorter100|2119_ ;
  assign \new_Sorter100|2220_  = \new_Sorter100|2120_  & \new_Sorter100|2121_ ;
  assign \new_Sorter100|2221_  = \new_Sorter100|2120_  | \new_Sorter100|2121_ ;
  assign \new_Sorter100|2222_  = \new_Sorter100|2122_  & \new_Sorter100|2123_ ;
  assign \new_Sorter100|2223_  = \new_Sorter100|2122_  | \new_Sorter100|2123_ ;
  assign \new_Sorter100|2224_  = \new_Sorter100|2124_  & \new_Sorter100|2125_ ;
  assign \new_Sorter100|2225_  = \new_Sorter100|2124_  | \new_Sorter100|2125_ ;
  assign \new_Sorter100|2226_  = \new_Sorter100|2126_  & \new_Sorter100|2127_ ;
  assign \new_Sorter100|2227_  = \new_Sorter100|2126_  | \new_Sorter100|2127_ ;
  assign \new_Sorter100|2228_  = \new_Sorter100|2128_  & \new_Sorter100|2129_ ;
  assign \new_Sorter100|2229_  = \new_Sorter100|2128_  | \new_Sorter100|2129_ ;
  assign \new_Sorter100|2230_  = \new_Sorter100|2130_  & \new_Sorter100|2131_ ;
  assign \new_Sorter100|2231_  = \new_Sorter100|2130_  | \new_Sorter100|2131_ ;
  assign \new_Sorter100|2232_  = \new_Sorter100|2132_  & \new_Sorter100|2133_ ;
  assign \new_Sorter100|2233_  = \new_Sorter100|2132_  | \new_Sorter100|2133_ ;
  assign \new_Sorter100|2234_  = \new_Sorter100|2134_  & \new_Sorter100|2135_ ;
  assign \new_Sorter100|2235_  = \new_Sorter100|2134_  | \new_Sorter100|2135_ ;
  assign \new_Sorter100|2236_  = \new_Sorter100|2136_  & \new_Sorter100|2137_ ;
  assign \new_Sorter100|2237_  = \new_Sorter100|2136_  | \new_Sorter100|2137_ ;
  assign \new_Sorter100|2238_  = \new_Sorter100|2138_  & \new_Sorter100|2139_ ;
  assign \new_Sorter100|2239_  = \new_Sorter100|2138_  | \new_Sorter100|2139_ ;
  assign \new_Sorter100|2240_  = \new_Sorter100|2140_  & \new_Sorter100|2141_ ;
  assign \new_Sorter100|2241_  = \new_Sorter100|2140_  | \new_Sorter100|2141_ ;
  assign \new_Sorter100|2242_  = \new_Sorter100|2142_  & \new_Sorter100|2143_ ;
  assign \new_Sorter100|2243_  = \new_Sorter100|2142_  | \new_Sorter100|2143_ ;
  assign \new_Sorter100|2244_  = \new_Sorter100|2144_  & \new_Sorter100|2145_ ;
  assign \new_Sorter100|2245_  = \new_Sorter100|2144_  | \new_Sorter100|2145_ ;
  assign \new_Sorter100|2246_  = \new_Sorter100|2146_  & \new_Sorter100|2147_ ;
  assign \new_Sorter100|2247_  = \new_Sorter100|2146_  | \new_Sorter100|2147_ ;
  assign \new_Sorter100|2248_  = \new_Sorter100|2148_  & \new_Sorter100|2149_ ;
  assign \new_Sorter100|2249_  = \new_Sorter100|2148_  | \new_Sorter100|2149_ ;
  assign \new_Sorter100|2250_  = \new_Sorter100|2150_  & \new_Sorter100|2151_ ;
  assign \new_Sorter100|2251_  = \new_Sorter100|2150_  | \new_Sorter100|2151_ ;
  assign \new_Sorter100|2252_  = \new_Sorter100|2152_  & \new_Sorter100|2153_ ;
  assign \new_Sorter100|2253_  = \new_Sorter100|2152_  | \new_Sorter100|2153_ ;
  assign \new_Sorter100|2254_  = \new_Sorter100|2154_  & \new_Sorter100|2155_ ;
  assign \new_Sorter100|2255_  = \new_Sorter100|2154_  | \new_Sorter100|2155_ ;
  assign \new_Sorter100|2256_  = \new_Sorter100|2156_  & \new_Sorter100|2157_ ;
  assign \new_Sorter100|2257_  = \new_Sorter100|2156_  | \new_Sorter100|2157_ ;
  assign \new_Sorter100|2258_  = \new_Sorter100|2158_  & \new_Sorter100|2159_ ;
  assign \new_Sorter100|2259_  = \new_Sorter100|2158_  | \new_Sorter100|2159_ ;
  assign \new_Sorter100|2260_  = \new_Sorter100|2160_  & \new_Sorter100|2161_ ;
  assign \new_Sorter100|2261_  = \new_Sorter100|2160_  | \new_Sorter100|2161_ ;
  assign \new_Sorter100|2262_  = \new_Sorter100|2162_  & \new_Sorter100|2163_ ;
  assign \new_Sorter100|2263_  = \new_Sorter100|2162_  | \new_Sorter100|2163_ ;
  assign \new_Sorter100|2264_  = \new_Sorter100|2164_  & \new_Sorter100|2165_ ;
  assign \new_Sorter100|2265_  = \new_Sorter100|2164_  | \new_Sorter100|2165_ ;
  assign \new_Sorter100|2266_  = \new_Sorter100|2166_  & \new_Sorter100|2167_ ;
  assign \new_Sorter100|2267_  = \new_Sorter100|2166_  | \new_Sorter100|2167_ ;
  assign \new_Sorter100|2268_  = \new_Sorter100|2168_  & \new_Sorter100|2169_ ;
  assign \new_Sorter100|2269_  = \new_Sorter100|2168_  | \new_Sorter100|2169_ ;
  assign \new_Sorter100|2270_  = \new_Sorter100|2170_  & \new_Sorter100|2171_ ;
  assign \new_Sorter100|2271_  = \new_Sorter100|2170_  | \new_Sorter100|2171_ ;
  assign \new_Sorter100|2272_  = \new_Sorter100|2172_  & \new_Sorter100|2173_ ;
  assign \new_Sorter100|2273_  = \new_Sorter100|2172_  | \new_Sorter100|2173_ ;
  assign \new_Sorter100|2274_  = \new_Sorter100|2174_  & \new_Sorter100|2175_ ;
  assign \new_Sorter100|2275_  = \new_Sorter100|2174_  | \new_Sorter100|2175_ ;
  assign \new_Sorter100|2276_  = \new_Sorter100|2176_  & \new_Sorter100|2177_ ;
  assign \new_Sorter100|2277_  = \new_Sorter100|2176_  | \new_Sorter100|2177_ ;
  assign \new_Sorter100|2278_  = \new_Sorter100|2178_  & \new_Sorter100|2179_ ;
  assign \new_Sorter100|2279_  = \new_Sorter100|2178_  | \new_Sorter100|2179_ ;
  assign \new_Sorter100|2280_  = \new_Sorter100|2180_  & \new_Sorter100|2181_ ;
  assign \new_Sorter100|2281_  = \new_Sorter100|2180_  | \new_Sorter100|2181_ ;
  assign \new_Sorter100|2282_  = \new_Sorter100|2182_  & \new_Sorter100|2183_ ;
  assign \new_Sorter100|2283_  = \new_Sorter100|2182_  | \new_Sorter100|2183_ ;
  assign \new_Sorter100|2284_  = \new_Sorter100|2184_  & \new_Sorter100|2185_ ;
  assign \new_Sorter100|2285_  = \new_Sorter100|2184_  | \new_Sorter100|2185_ ;
  assign \new_Sorter100|2286_  = \new_Sorter100|2186_  & \new_Sorter100|2187_ ;
  assign \new_Sorter100|2287_  = \new_Sorter100|2186_  | \new_Sorter100|2187_ ;
  assign \new_Sorter100|2288_  = \new_Sorter100|2188_  & \new_Sorter100|2189_ ;
  assign \new_Sorter100|2289_  = \new_Sorter100|2188_  | \new_Sorter100|2189_ ;
  assign \new_Sorter100|2290_  = \new_Sorter100|2190_  & \new_Sorter100|2191_ ;
  assign \new_Sorter100|2291_  = \new_Sorter100|2190_  | \new_Sorter100|2191_ ;
  assign \new_Sorter100|2292_  = \new_Sorter100|2192_  & \new_Sorter100|2193_ ;
  assign \new_Sorter100|2293_  = \new_Sorter100|2192_  | \new_Sorter100|2193_ ;
  assign \new_Sorter100|2294_  = \new_Sorter100|2194_  & \new_Sorter100|2195_ ;
  assign \new_Sorter100|2295_  = \new_Sorter100|2194_  | \new_Sorter100|2195_ ;
  assign \new_Sorter100|2296_  = \new_Sorter100|2196_  & \new_Sorter100|2197_ ;
  assign \new_Sorter100|2297_  = \new_Sorter100|2196_  | \new_Sorter100|2197_ ;
  assign \new_Sorter100|2298_  = \new_Sorter100|2198_  & \new_Sorter100|2199_ ;
  assign \new_Sorter100|2299_  = \new_Sorter100|2198_  | \new_Sorter100|2199_ ;
  assign \new_Sorter100|2300_  = \new_Sorter100|2200_ ;
  assign \new_Sorter100|2399_  = \new_Sorter100|2299_ ;
  assign \new_Sorter100|2301_  = \new_Sorter100|2201_  & \new_Sorter100|2202_ ;
  assign \new_Sorter100|2302_  = \new_Sorter100|2201_  | \new_Sorter100|2202_ ;
  assign \new_Sorter100|2303_  = \new_Sorter100|2203_  & \new_Sorter100|2204_ ;
  assign \new_Sorter100|2304_  = \new_Sorter100|2203_  | \new_Sorter100|2204_ ;
  assign \new_Sorter100|2305_  = \new_Sorter100|2205_  & \new_Sorter100|2206_ ;
  assign \new_Sorter100|2306_  = \new_Sorter100|2205_  | \new_Sorter100|2206_ ;
  assign \new_Sorter100|2307_  = \new_Sorter100|2207_  & \new_Sorter100|2208_ ;
  assign \new_Sorter100|2308_  = \new_Sorter100|2207_  | \new_Sorter100|2208_ ;
  assign \new_Sorter100|2309_  = \new_Sorter100|2209_  & \new_Sorter100|2210_ ;
  assign \new_Sorter100|2310_  = \new_Sorter100|2209_  | \new_Sorter100|2210_ ;
  assign \new_Sorter100|2311_  = \new_Sorter100|2211_  & \new_Sorter100|2212_ ;
  assign \new_Sorter100|2312_  = \new_Sorter100|2211_  | \new_Sorter100|2212_ ;
  assign \new_Sorter100|2313_  = \new_Sorter100|2213_  & \new_Sorter100|2214_ ;
  assign \new_Sorter100|2314_  = \new_Sorter100|2213_  | \new_Sorter100|2214_ ;
  assign \new_Sorter100|2315_  = \new_Sorter100|2215_  & \new_Sorter100|2216_ ;
  assign \new_Sorter100|2316_  = \new_Sorter100|2215_  | \new_Sorter100|2216_ ;
  assign \new_Sorter100|2317_  = \new_Sorter100|2217_  & \new_Sorter100|2218_ ;
  assign \new_Sorter100|2318_  = \new_Sorter100|2217_  | \new_Sorter100|2218_ ;
  assign \new_Sorter100|2319_  = \new_Sorter100|2219_  & \new_Sorter100|2220_ ;
  assign \new_Sorter100|2320_  = \new_Sorter100|2219_  | \new_Sorter100|2220_ ;
  assign \new_Sorter100|2321_  = \new_Sorter100|2221_  & \new_Sorter100|2222_ ;
  assign \new_Sorter100|2322_  = \new_Sorter100|2221_  | \new_Sorter100|2222_ ;
  assign \new_Sorter100|2323_  = \new_Sorter100|2223_  & \new_Sorter100|2224_ ;
  assign \new_Sorter100|2324_  = \new_Sorter100|2223_  | \new_Sorter100|2224_ ;
  assign \new_Sorter100|2325_  = \new_Sorter100|2225_  & \new_Sorter100|2226_ ;
  assign \new_Sorter100|2326_  = \new_Sorter100|2225_  | \new_Sorter100|2226_ ;
  assign \new_Sorter100|2327_  = \new_Sorter100|2227_  & \new_Sorter100|2228_ ;
  assign \new_Sorter100|2328_  = \new_Sorter100|2227_  | \new_Sorter100|2228_ ;
  assign \new_Sorter100|2329_  = \new_Sorter100|2229_  & \new_Sorter100|2230_ ;
  assign \new_Sorter100|2330_  = \new_Sorter100|2229_  | \new_Sorter100|2230_ ;
  assign \new_Sorter100|2331_  = \new_Sorter100|2231_  & \new_Sorter100|2232_ ;
  assign \new_Sorter100|2332_  = \new_Sorter100|2231_  | \new_Sorter100|2232_ ;
  assign \new_Sorter100|2333_  = \new_Sorter100|2233_  & \new_Sorter100|2234_ ;
  assign \new_Sorter100|2334_  = \new_Sorter100|2233_  | \new_Sorter100|2234_ ;
  assign \new_Sorter100|2335_  = \new_Sorter100|2235_  & \new_Sorter100|2236_ ;
  assign \new_Sorter100|2336_  = \new_Sorter100|2235_  | \new_Sorter100|2236_ ;
  assign \new_Sorter100|2337_  = \new_Sorter100|2237_  & \new_Sorter100|2238_ ;
  assign \new_Sorter100|2338_  = \new_Sorter100|2237_  | \new_Sorter100|2238_ ;
  assign \new_Sorter100|2339_  = \new_Sorter100|2239_  & \new_Sorter100|2240_ ;
  assign \new_Sorter100|2340_  = \new_Sorter100|2239_  | \new_Sorter100|2240_ ;
  assign \new_Sorter100|2341_  = \new_Sorter100|2241_  & \new_Sorter100|2242_ ;
  assign \new_Sorter100|2342_  = \new_Sorter100|2241_  | \new_Sorter100|2242_ ;
  assign \new_Sorter100|2343_  = \new_Sorter100|2243_  & \new_Sorter100|2244_ ;
  assign \new_Sorter100|2344_  = \new_Sorter100|2243_  | \new_Sorter100|2244_ ;
  assign \new_Sorter100|2345_  = \new_Sorter100|2245_  & \new_Sorter100|2246_ ;
  assign \new_Sorter100|2346_  = \new_Sorter100|2245_  | \new_Sorter100|2246_ ;
  assign \new_Sorter100|2347_  = \new_Sorter100|2247_  & \new_Sorter100|2248_ ;
  assign \new_Sorter100|2348_  = \new_Sorter100|2247_  | \new_Sorter100|2248_ ;
  assign \new_Sorter100|2349_  = \new_Sorter100|2249_  & \new_Sorter100|2250_ ;
  assign \new_Sorter100|2350_  = \new_Sorter100|2249_  | \new_Sorter100|2250_ ;
  assign \new_Sorter100|2351_  = \new_Sorter100|2251_  & \new_Sorter100|2252_ ;
  assign \new_Sorter100|2352_  = \new_Sorter100|2251_  | \new_Sorter100|2252_ ;
  assign \new_Sorter100|2353_  = \new_Sorter100|2253_  & \new_Sorter100|2254_ ;
  assign \new_Sorter100|2354_  = \new_Sorter100|2253_  | \new_Sorter100|2254_ ;
  assign \new_Sorter100|2355_  = \new_Sorter100|2255_  & \new_Sorter100|2256_ ;
  assign \new_Sorter100|2356_  = \new_Sorter100|2255_  | \new_Sorter100|2256_ ;
  assign \new_Sorter100|2357_  = \new_Sorter100|2257_  & \new_Sorter100|2258_ ;
  assign \new_Sorter100|2358_  = \new_Sorter100|2257_  | \new_Sorter100|2258_ ;
  assign \new_Sorter100|2359_  = \new_Sorter100|2259_  & \new_Sorter100|2260_ ;
  assign \new_Sorter100|2360_  = \new_Sorter100|2259_  | \new_Sorter100|2260_ ;
  assign \new_Sorter100|2361_  = \new_Sorter100|2261_  & \new_Sorter100|2262_ ;
  assign \new_Sorter100|2362_  = \new_Sorter100|2261_  | \new_Sorter100|2262_ ;
  assign \new_Sorter100|2363_  = \new_Sorter100|2263_  & \new_Sorter100|2264_ ;
  assign \new_Sorter100|2364_  = \new_Sorter100|2263_  | \new_Sorter100|2264_ ;
  assign \new_Sorter100|2365_  = \new_Sorter100|2265_  & \new_Sorter100|2266_ ;
  assign \new_Sorter100|2366_  = \new_Sorter100|2265_  | \new_Sorter100|2266_ ;
  assign \new_Sorter100|2367_  = \new_Sorter100|2267_  & \new_Sorter100|2268_ ;
  assign \new_Sorter100|2368_  = \new_Sorter100|2267_  | \new_Sorter100|2268_ ;
  assign \new_Sorter100|2369_  = \new_Sorter100|2269_  & \new_Sorter100|2270_ ;
  assign \new_Sorter100|2370_  = \new_Sorter100|2269_  | \new_Sorter100|2270_ ;
  assign \new_Sorter100|2371_  = \new_Sorter100|2271_  & \new_Sorter100|2272_ ;
  assign \new_Sorter100|2372_  = \new_Sorter100|2271_  | \new_Sorter100|2272_ ;
  assign \new_Sorter100|2373_  = \new_Sorter100|2273_  & \new_Sorter100|2274_ ;
  assign \new_Sorter100|2374_  = \new_Sorter100|2273_  | \new_Sorter100|2274_ ;
  assign \new_Sorter100|2375_  = \new_Sorter100|2275_  & \new_Sorter100|2276_ ;
  assign \new_Sorter100|2376_  = \new_Sorter100|2275_  | \new_Sorter100|2276_ ;
  assign \new_Sorter100|2377_  = \new_Sorter100|2277_  & \new_Sorter100|2278_ ;
  assign \new_Sorter100|2378_  = \new_Sorter100|2277_  | \new_Sorter100|2278_ ;
  assign \new_Sorter100|2379_  = \new_Sorter100|2279_  & \new_Sorter100|2280_ ;
  assign \new_Sorter100|2380_  = \new_Sorter100|2279_  | \new_Sorter100|2280_ ;
  assign \new_Sorter100|2381_  = \new_Sorter100|2281_  & \new_Sorter100|2282_ ;
  assign \new_Sorter100|2382_  = \new_Sorter100|2281_  | \new_Sorter100|2282_ ;
  assign \new_Sorter100|2383_  = \new_Sorter100|2283_  & \new_Sorter100|2284_ ;
  assign \new_Sorter100|2384_  = \new_Sorter100|2283_  | \new_Sorter100|2284_ ;
  assign \new_Sorter100|2385_  = \new_Sorter100|2285_  & \new_Sorter100|2286_ ;
  assign \new_Sorter100|2386_  = \new_Sorter100|2285_  | \new_Sorter100|2286_ ;
  assign \new_Sorter100|2387_  = \new_Sorter100|2287_  & \new_Sorter100|2288_ ;
  assign \new_Sorter100|2388_  = \new_Sorter100|2287_  | \new_Sorter100|2288_ ;
  assign \new_Sorter100|2389_  = \new_Sorter100|2289_  & \new_Sorter100|2290_ ;
  assign \new_Sorter100|2390_  = \new_Sorter100|2289_  | \new_Sorter100|2290_ ;
  assign \new_Sorter100|2391_  = \new_Sorter100|2291_  & \new_Sorter100|2292_ ;
  assign \new_Sorter100|2392_  = \new_Sorter100|2291_  | \new_Sorter100|2292_ ;
  assign \new_Sorter100|2393_  = \new_Sorter100|2293_  & \new_Sorter100|2294_ ;
  assign \new_Sorter100|2394_  = \new_Sorter100|2293_  | \new_Sorter100|2294_ ;
  assign \new_Sorter100|2395_  = \new_Sorter100|2295_  & \new_Sorter100|2296_ ;
  assign \new_Sorter100|2396_  = \new_Sorter100|2295_  | \new_Sorter100|2296_ ;
  assign \new_Sorter100|2397_  = \new_Sorter100|2297_  & \new_Sorter100|2298_ ;
  assign \new_Sorter100|2398_  = \new_Sorter100|2297_  | \new_Sorter100|2298_ ;
  assign \new_Sorter100|2400_  = \new_Sorter100|2300_  & \new_Sorter100|2301_ ;
  assign \new_Sorter100|2401_  = \new_Sorter100|2300_  | \new_Sorter100|2301_ ;
  assign \new_Sorter100|2402_  = \new_Sorter100|2302_  & \new_Sorter100|2303_ ;
  assign \new_Sorter100|2403_  = \new_Sorter100|2302_  | \new_Sorter100|2303_ ;
  assign \new_Sorter100|2404_  = \new_Sorter100|2304_  & \new_Sorter100|2305_ ;
  assign \new_Sorter100|2405_  = \new_Sorter100|2304_  | \new_Sorter100|2305_ ;
  assign \new_Sorter100|2406_  = \new_Sorter100|2306_  & \new_Sorter100|2307_ ;
  assign \new_Sorter100|2407_  = \new_Sorter100|2306_  | \new_Sorter100|2307_ ;
  assign \new_Sorter100|2408_  = \new_Sorter100|2308_  & \new_Sorter100|2309_ ;
  assign \new_Sorter100|2409_  = \new_Sorter100|2308_  | \new_Sorter100|2309_ ;
  assign \new_Sorter100|2410_  = \new_Sorter100|2310_  & \new_Sorter100|2311_ ;
  assign \new_Sorter100|2411_  = \new_Sorter100|2310_  | \new_Sorter100|2311_ ;
  assign \new_Sorter100|2412_  = \new_Sorter100|2312_  & \new_Sorter100|2313_ ;
  assign \new_Sorter100|2413_  = \new_Sorter100|2312_  | \new_Sorter100|2313_ ;
  assign \new_Sorter100|2414_  = \new_Sorter100|2314_  & \new_Sorter100|2315_ ;
  assign \new_Sorter100|2415_  = \new_Sorter100|2314_  | \new_Sorter100|2315_ ;
  assign \new_Sorter100|2416_  = \new_Sorter100|2316_  & \new_Sorter100|2317_ ;
  assign \new_Sorter100|2417_  = \new_Sorter100|2316_  | \new_Sorter100|2317_ ;
  assign \new_Sorter100|2418_  = \new_Sorter100|2318_  & \new_Sorter100|2319_ ;
  assign \new_Sorter100|2419_  = \new_Sorter100|2318_  | \new_Sorter100|2319_ ;
  assign \new_Sorter100|2420_  = \new_Sorter100|2320_  & \new_Sorter100|2321_ ;
  assign \new_Sorter100|2421_  = \new_Sorter100|2320_  | \new_Sorter100|2321_ ;
  assign \new_Sorter100|2422_  = \new_Sorter100|2322_  & \new_Sorter100|2323_ ;
  assign \new_Sorter100|2423_  = \new_Sorter100|2322_  | \new_Sorter100|2323_ ;
  assign \new_Sorter100|2424_  = \new_Sorter100|2324_  & \new_Sorter100|2325_ ;
  assign \new_Sorter100|2425_  = \new_Sorter100|2324_  | \new_Sorter100|2325_ ;
  assign \new_Sorter100|2426_  = \new_Sorter100|2326_  & \new_Sorter100|2327_ ;
  assign \new_Sorter100|2427_  = \new_Sorter100|2326_  | \new_Sorter100|2327_ ;
  assign \new_Sorter100|2428_  = \new_Sorter100|2328_  & \new_Sorter100|2329_ ;
  assign \new_Sorter100|2429_  = \new_Sorter100|2328_  | \new_Sorter100|2329_ ;
  assign \new_Sorter100|2430_  = \new_Sorter100|2330_  & \new_Sorter100|2331_ ;
  assign \new_Sorter100|2431_  = \new_Sorter100|2330_  | \new_Sorter100|2331_ ;
  assign \new_Sorter100|2432_  = \new_Sorter100|2332_  & \new_Sorter100|2333_ ;
  assign \new_Sorter100|2433_  = \new_Sorter100|2332_  | \new_Sorter100|2333_ ;
  assign \new_Sorter100|2434_  = \new_Sorter100|2334_  & \new_Sorter100|2335_ ;
  assign \new_Sorter100|2435_  = \new_Sorter100|2334_  | \new_Sorter100|2335_ ;
  assign \new_Sorter100|2436_  = \new_Sorter100|2336_  & \new_Sorter100|2337_ ;
  assign \new_Sorter100|2437_  = \new_Sorter100|2336_  | \new_Sorter100|2337_ ;
  assign \new_Sorter100|2438_  = \new_Sorter100|2338_  & \new_Sorter100|2339_ ;
  assign \new_Sorter100|2439_  = \new_Sorter100|2338_  | \new_Sorter100|2339_ ;
  assign \new_Sorter100|2440_  = \new_Sorter100|2340_  & \new_Sorter100|2341_ ;
  assign \new_Sorter100|2441_  = \new_Sorter100|2340_  | \new_Sorter100|2341_ ;
  assign \new_Sorter100|2442_  = \new_Sorter100|2342_  & \new_Sorter100|2343_ ;
  assign \new_Sorter100|2443_  = \new_Sorter100|2342_  | \new_Sorter100|2343_ ;
  assign \new_Sorter100|2444_  = \new_Sorter100|2344_  & \new_Sorter100|2345_ ;
  assign \new_Sorter100|2445_  = \new_Sorter100|2344_  | \new_Sorter100|2345_ ;
  assign \new_Sorter100|2446_  = \new_Sorter100|2346_  & \new_Sorter100|2347_ ;
  assign \new_Sorter100|2447_  = \new_Sorter100|2346_  | \new_Sorter100|2347_ ;
  assign \new_Sorter100|2448_  = \new_Sorter100|2348_  & \new_Sorter100|2349_ ;
  assign \new_Sorter100|2449_  = \new_Sorter100|2348_  | \new_Sorter100|2349_ ;
  assign \new_Sorter100|2450_  = \new_Sorter100|2350_  & \new_Sorter100|2351_ ;
  assign \new_Sorter100|2451_  = \new_Sorter100|2350_  | \new_Sorter100|2351_ ;
  assign \new_Sorter100|2452_  = \new_Sorter100|2352_  & \new_Sorter100|2353_ ;
  assign \new_Sorter100|2453_  = \new_Sorter100|2352_  | \new_Sorter100|2353_ ;
  assign \new_Sorter100|2454_  = \new_Sorter100|2354_  & \new_Sorter100|2355_ ;
  assign \new_Sorter100|2455_  = \new_Sorter100|2354_  | \new_Sorter100|2355_ ;
  assign \new_Sorter100|2456_  = \new_Sorter100|2356_  & \new_Sorter100|2357_ ;
  assign \new_Sorter100|2457_  = \new_Sorter100|2356_  | \new_Sorter100|2357_ ;
  assign \new_Sorter100|2458_  = \new_Sorter100|2358_  & \new_Sorter100|2359_ ;
  assign \new_Sorter100|2459_  = \new_Sorter100|2358_  | \new_Sorter100|2359_ ;
  assign \new_Sorter100|2460_  = \new_Sorter100|2360_  & \new_Sorter100|2361_ ;
  assign \new_Sorter100|2461_  = \new_Sorter100|2360_  | \new_Sorter100|2361_ ;
  assign \new_Sorter100|2462_  = \new_Sorter100|2362_  & \new_Sorter100|2363_ ;
  assign \new_Sorter100|2463_  = \new_Sorter100|2362_  | \new_Sorter100|2363_ ;
  assign \new_Sorter100|2464_  = \new_Sorter100|2364_  & \new_Sorter100|2365_ ;
  assign \new_Sorter100|2465_  = \new_Sorter100|2364_  | \new_Sorter100|2365_ ;
  assign \new_Sorter100|2466_  = \new_Sorter100|2366_  & \new_Sorter100|2367_ ;
  assign \new_Sorter100|2467_  = \new_Sorter100|2366_  | \new_Sorter100|2367_ ;
  assign \new_Sorter100|2468_  = \new_Sorter100|2368_  & \new_Sorter100|2369_ ;
  assign \new_Sorter100|2469_  = \new_Sorter100|2368_  | \new_Sorter100|2369_ ;
  assign \new_Sorter100|2470_  = \new_Sorter100|2370_  & \new_Sorter100|2371_ ;
  assign \new_Sorter100|2471_  = \new_Sorter100|2370_  | \new_Sorter100|2371_ ;
  assign \new_Sorter100|2472_  = \new_Sorter100|2372_  & \new_Sorter100|2373_ ;
  assign \new_Sorter100|2473_  = \new_Sorter100|2372_  | \new_Sorter100|2373_ ;
  assign \new_Sorter100|2474_  = \new_Sorter100|2374_  & \new_Sorter100|2375_ ;
  assign \new_Sorter100|2475_  = \new_Sorter100|2374_  | \new_Sorter100|2375_ ;
  assign \new_Sorter100|2476_  = \new_Sorter100|2376_  & \new_Sorter100|2377_ ;
  assign \new_Sorter100|2477_  = \new_Sorter100|2376_  | \new_Sorter100|2377_ ;
  assign \new_Sorter100|2478_  = \new_Sorter100|2378_  & \new_Sorter100|2379_ ;
  assign \new_Sorter100|2479_  = \new_Sorter100|2378_  | \new_Sorter100|2379_ ;
  assign \new_Sorter100|2480_  = \new_Sorter100|2380_  & \new_Sorter100|2381_ ;
  assign \new_Sorter100|2481_  = \new_Sorter100|2380_  | \new_Sorter100|2381_ ;
  assign \new_Sorter100|2482_  = \new_Sorter100|2382_  & \new_Sorter100|2383_ ;
  assign \new_Sorter100|2483_  = \new_Sorter100|2382_  | \new_Sorter100|2383_ ;
  assign \new_Sorter100|2484_  = \new_Sorter100|2384_  & \new_Sorter100|2385_ ;
  assign \new_Sorter100|2485_  = \new_Sorter100|2384_  | \new_Sorter100|2385_ ;
  assign \new_Sorter100|2486_  = \new_Sorter100|2386_  & \new_Sorter100|2387_ ;
  assign \new_Sorter100|2487_  = \new_Sorter100|2386_  | \new_Sorter100|2387_ ;
  assign \new_Sorter100|2488_  = \new_Sorter100|2388_  & \new_Sorter100|2389_ ;
  assign \new_Sorter100|2489_  = \new_Sorter100|2388_  | \new_Sorter100|2389_ ;
  assign \new_Sorter100|2490_  = \new_Sorter100|2390_  & \new_Sorter100|2391_ ;
  assign \new_Sorter100|2491_  = \new_Sorter100|2390_  | \new_Sorter100|2391_ ;
  assign \new_Sorter100|2492_  = \new_Sorter100|2392_  & \new_Sorter100|2393_ ;
  assign \new_Sorter100|2493_  = \new_Sorter100|2392_  | \new_Sorter100|2393_ ;
  assign \new_Sorter100|2494_  = \new_Sorter100|2394_  & \new_Sorter100|2395_ ;
  assign \new_Sorter100|2495_  = \new_Sorter100|2394_  | \new_Sorter100|2395_ ;
  assign \new_Sorter100|2496_  = \new_Sorter100|2396_  & \new_Sorter100|2397_ ;
  assign \new_Sorter100|2497_  = \new_Sorter100|2396_  | \new_Sorter100|2397_ ;
  assign \new_Sorter100|2498_  = \new_Sorter100|2398_  & \new_Sorter100|2399_ ;
  assign \new_Sorter100|2499_  = \new_Sorter100|2398_  | \new_Sorter100|2399_ ;
  assign \new_Sorter100|2500_  = \new_Sorter100|2400_ ;
  assign \new_Sorter100|2599_  = \new_Sorter100|2499_ ;
  assign \new_Sorter100|2501_  = \new_Sorter100|2401_  & \new_Sorter100|2402_ ;
  assign \new_Sorter100|2502_  = \new_Sorter100|2401_  | \new_Sorter100|2402_ ;
  assign \new_Sorter100|2503_  = \new_Sorter100|2403_  & \new_Sorter100|2404_ ;
  assign \new_Sorter100|2504_  = \new_Sorter100|2403_  | \new_Sorter100|2404_ ;
  assign \new_Sorter100|2505_  = \new_Sorter100|2405_  & \new_Sorter100|2406_ ;
  assign \new_Sorter100|2506_  = \new_Sorter100|2405_  | \new_Sorter100|2406_ ;
  assign \new_Sorter100|2507_  = \new_Sorter100|2407_  & \new_Sorter100|2408_ ;
  assign \new_Sorter100|2508_  = \new_Sorter100|2407_  | \new_Sorter100|2408_ ;
  assign \new_Sorter100|2509_  = \new_Sorter100|2409_  & \new_Sorter100|2410_ ;
  assign \new_Sorter100|2510_  = \new_Sorter100|2409_  | \new_Sorter100|2410_ ;
  assign \new_Sorter100|2511_  = \new_Sorter100|2411_  & \new_Sorter100|2412_ ;
  assign \new_Sorter100|2512_  = \new_Sorter100|2411_  | \new_Sorter100|2412_ ;
  assign \new_Sorter100|2513_  = \new_Sorter100|2413_  & \new_Sorter100|2414_ ;
  assign \new_Sorter100|2514_  = \new_Sorter100|2413_  | \new_Sorter100|2414_ ;
  assign \new_Sorter100|2515_  = \new_Sorter100|2415_  & \new_Sorter100|2416_ ;
  assign \new_Sorter100|2516_  = \new_Sorter100|2415_  | \new_Sorter100|2416_ ;
  assign \new_Sorter100|2517_  = \new_Sorter100|2417_  & \new_Sorter100|2418_ ;
  assign \new_Sorter100|2518_  = \new_Sorter100|2417_  | \new_Sorter100|2418_ ;
  assign \new_Sorter100|2519_  = \new_Sorter100|2419_  & \new_Sorter100|2420_ ;
  assign \new_Sorter100|2520_  = \new_Sorter100|2419_  | \new_Sorter100|2420_ ;
  assign \new_Sorter100|2521_  = \new_Sorter100|2421_  & \new_Sorter100|2422_ ;
  assign \new_Sorter100|2522_  = \new_Sorter100|2421_  | \new_Sorter100|2422_ ;
  assign \new_Sorter100|2523_  = \new_Sorter100|2423_  & \new_Sorter100|2424_ ;
  assign \new_Sorter100|2524_  = \new_Sorter100|2423_  | \new_Sorter100|2424_ ;
  assign \new_Sorter100|2525_  = \new_Sorter100|2425_  & \new_Sorter100|2426_ ;
  assign \new_Sorter100|2526_  = \new_Sorter100|2425_  | \new_Sorter100|2426_ ;
  assign \new_Sorter100|2527_  = \new_Sorter100|2427_  & \new_Sorter100|2428_ ;
  assign \new_Sorter100|2528_  = \new_Sorter100|2427_  | \new_Sorter100|2428_ ;
  assign \new_Sorter100|2529_  = \new_Sorter100|2429_  & \new_Sorter100|2430_ ;
  assign \new_Sorter100|2530_  = \new_Sorter100|2429_  | \new_Sorter100|2430_ ;
  assign \new_Sorter100|2531_  = \new_Sorter100|2431_  & \new_Sorter100|2432_ ;
  assign \new_Sorter100|2532_  = \new_Sorter100|2431_  | \new_Sorter100|2432_ ;
  assign \new_Sorter100|2533_  = \new_Sorter100|2433_  & \new_Sorter100|2434_ ;
  assign \new_Sorter100|2534_  = \new_Sorter100|2433_  | \new_Sorter100|2434_ ;
  assign \new_Sorter100|2535_  = \new_Sorter100|2435_  & \new_Sorter100|2436_ ;
  assign \new_Sorter100|2536_  = \new_Sorter100|2435_  | \new_Sorter100|2436_ ;
  assign \new_Sorter100|2537_  = \new_Sorter100|2437_  & \new_Sorter100|2438_ ;
  assign \new_Sorter100|2538_  = \new_Sorter100|2437_  | \new_Sorter100|2438_ ;
  assign \new_Sorter100|2539_  = \new_Sorter100|2439_  & \new_Sorter100|2440_ ;
  assign \new_Sorter100|2540_  = \new_Sorter100|2439_  | \new_Sorter100|2440_ ;
  assign \new_Sorter100|2541_  = \new_Sorter100|2441_  & \new_Sorter100|2442_ ;
  assign \new_Sorter100|2542_  = \new_Sorter100|2441_  | \new_Sorter100|2442_ ;
  assign \new_Sorter100|2543_  = \new_Sorter100|2443_  & \new_Sorter100|2444_ ;
  assign \new_Sorter100|2544_  = \new_Sorter100|2443_  | \new_Sorter100|2444_ ;
  assign \new_Sorter100|2545_  = \new_Sorter100|2445_  & \new_Sorter100|2446_ ;
  assign \new_Sorter100|2546_  = \new_Sorter100|2445_  | \new_Sorter100|2446_ ;
  assign \new_Sorter100|2547_  = \new_Sorter100|2447_  & \new_Sorter100|2448_ ;
  assign \new_Sorter100|2548_  = \new_Sorter100|2447_  | \new_Sorter100|2448_ ;
  assign \new_Sorter100|2549_  = \new_Sorter100|2449_  & \new_Sorter100|2450_ ;
  assign \new_Sorter100|2550_  = \new_Sorter100|2449_  | \new_Sorter100|2450_ ;
  assign \new_Sorter100|2551_  = \new_Sorter100|2451_  & \new_Sorter100|2452_ ;
  assign \new_Sorter100|2552_  = \new_Sorter100|2451_  | \new_Sorter100|2452_ ;
  assign \new_Sorter100|2553_  = \new_Sorter100|2453_  & \new_Sorter100|2454_ ;
  assign \new_Sorter100|2554_  = \new_Sorter100|2453_  | \new_Sorter100|2454_ ;
  assign \new_Sorter100|2555_  = \new_Sorter100|2455_  & \new_Sorter100|2456_ ;
  assign \new_Sorter100|2556_  = \new_Sorter100|2455_  | \new_Sorter100|2456_ ;
  assign \new_Sorter100|2557_  = \new_Sorter100|2457_  & \new_Sorter100|2458_ ;
  assign \new_Sorter100|2558_  = \new_Sorter100|2457_  | \new_Sorter100|2458_ ;
  assign \new_Sorter100|2559_  = \new_Sorter100|2459_  & \new_Sorter100|2460_ ;
  assign \new_Sorter100|2560_  = \new_Sorter100|2459_  | \new_Sorter100|2460_ ;
  assign \new_Sorter100|2561_  = \new_Sorter100|2461_  & \new_Sorter100|2462_ ;
  assign \new_Sorter100|2562_  = \new_Sorter100|2461_  | \new_Sorter100|2462_ ;
  assign \new_Sorter100|2563_  = \new_Sorter100|2463_  & \new_Sorter100|2464_ ;
  assign \new_Sorter100|2564_  = \new_Sorter100|2463_  | \new_Sorter100|2464_ ;
  assign \new_Sorter100|2565_  = \new_Sorter100|2465_  & \new_Sorter100|2466_ ;
  assign \new_Sorter100|2566_  = \new_Sorter100|2465_  | \new_Sorter100|2466_ ;
  assign \new_Sorter100|2567_  = \new_Sorter100|2467_  & \new_Sorter100|2468_ ;
  assign \new_Sorter100|2568_  = \new_Sorter100|2467_  | \new_Sorter100|2468_ ;
  assign \new_Sorter100|2569_  = \new_Sorter100|2469_  & \new_Sorter100|2470_ ;
  assign \new_Sorter100|2570_  = \new_Sorter100|2469_  | \new_Sorter100|2470_ ;
  assign \new_Sorter100|2571_  = \new_Sorter100|2471_  & \new_Sorter100|2472_ ;
  assign \new_Sorter100|2572_  = \new_Sorter100|2471_  | \new_Sorter100|2472_ ;
  assign \new_Sorter100|2573_  = \new_Sorter100|2473_  & \new_Sorter100|2474_ ;
  assign \new_Sorter100|2574_  = \new_Sorter100|2473_  | \new_Sorter100|2474_ ;
  assign \new_Sorter100|2575_  = \new_Sorter100|2475_  & \new_Sorter100|2476_ ;
  assign \new_Sorter100|2576_  = \new_Sorter100|2475_  | \new_Sorter100|2476_ ;
  assign \new_Sorter100|2577_  = \new_Sorter100|2477_  & \new_Sorter100|2478_ ;
  assign \new_Sorter100|2578_  = \new_Sorter100|2477_  | \new_Sorter100|2478_ ;
  assign \new_Sorter100|2579_  = \new_Sorter100|2479_  & \new_Sorter100|2480_ ;
  assign \new_Sorter100|2580_  = \new_Sorter100|2479_  | \new_Sorter100|2480_ ;
  assign \new_Sorter100|2581_  = \new_Sorter100|2481_  & \new_Sorter100|2482_ ;
  assign \new_Sorter100|2582_  = \new_Sorter100|2481_  | \new_Sorter100|2482_ ;
  assign \new_Sorter100|2583_  = \new_Sorter100|2483_  & \new_Sorter100|2484_ ;
  assign \new_Sorter100|2584_  = \new_Sorter100|2483_  | \new_Sorter100|2484_ ;
  assign \new_Sorter100|2585_  = \new_Sorter100|2485_  & \new_Sorter100|2486_ ;
  assign \new_Sorter100|2586_  = \new_Sorter100|2485_  | \new_Sorter100|2486_ ;
  assign \new_Sorter100|2587_  = \new_Sorter100|2487_  & \new_Sorter100|2488_ ;
  assign \new_Sorter100|2588_  = \new_Sorter100|2487_  | \new_Sorter100|2488_ ;
  assign \new_Sorter100|2589_  = \new_Sorter100|2489_  & \new_Sorter100|2490_ ;
  assign \new_Sorter100|2590_  = \new_Sorter100|2489_  | \new_Sorter100|2490_ ;
  assign \new_Sorter100|2591_  = \new_Sorter100|2491_  & \new_Sorter100|2492_ ;
  assign \new_Sorter100|2592_  = \new_Sorter100|2491_  | \new_Sorter100|2492_ ;
  assign \new_Sorter100|2593_  = \new_Sorter100|2493_  & \new_Sorter100|2494_ ;
  assign \new_Sorter100|2594_  = \new_Sorter100|2493_  | \new_Sorter100|2494_ ;
  assign \new_Sorter100|2595_  = \new_Sorter100|2495_  & \new_Sorter100|2496_ ;
  assign \new_Sorter100|2596_  = \new_Sorter100|2495_  | \new_Sorter100|2496_ ;
  assign \new_Sorter100|2597_  = \new_Sorter100|2497_  & \new_Sorter100|2498_ ;
  assign \new_Sorter100|2598_  = \new_Sorter100|2497_  | \new_Sorter100|2498_ ;
  assign \new_Sorter100|2600_  = \new_Sorter100|2500_  & \new_Sorter100|2501_ ;
  assign \new_Sorter100|2601_  = \new_Sorter100|2500_  | \new_Sorter100|2501_ ;
  assign \new_Sorter100|2602_  = \new_Sorter100|2502_  & \new_Sorter100|2503_ ;
  assign \new_Sorter100|2603_  = \new_Sorter100|2502_  | \new_Sorter100|2503_ ;
  assign \new_Sorter100|2604_  = \new_Sorter100|2504_  & \new_Sorter100|2505_ ;
  assign \new_Sorter100|2605_  = \new_Sorter100|2504_  | \new_Sorter100|2505_ ;
  assign \new_Sorter100|2606_  = \new_Sorter100|2506_  & \new_Sorter100|2507_ ;
  assign \new_Sorter100|2607_  = \new_Sorter100|2506_  | \new_Sorter100|2507_ ;
  assign \new_Sorter100|2608_  = \new_Sorter100|2508_  & \new_Sorter100|2509_ ;
  assign \new_Sorter100|2609_  = \new_Sorter100|2508_  | \new_Sorter100|2509_ ;
  assign \new_Sorter100|2610_  = \new_Sorter100|2510_  & \new_Sorter100|2511_ ;
  assign \new_Sorter100|2611_  = \new_Sorter100|2510_  | \new_Sorter100|2511_ ;
  assign \new_Sorter100|2612_  = \new_Sorter100|2512_  & \new_Sorter100|2513_ ;
  assign \new_Sorter100|2613_  = \new_Sorter100|2512_  | \new_Sorter100|2513_ ;
  assign \new_Sorter100|2614_  = \new_Sorter100|2514_  & \new_Sorter100|2515_ ;
  assign \new_Sorter100|2615_  = \new_Sorter100|2514_  | \new_Sorter100|2515_ ;
  assign \new_Sorter100|2616_  = \new_Sorter100|2516_  & \new_Sorter100|2517_ ;
  assign \new_Sorter100|2617_  = \new_Sorter100|2516_  | \new_Sorter100|2517_ ;
  assign \new_Sorter100|2618_  = \new_Sorter100|2518_  & \new_Sorter100|2519_ ;
  assign \new_Sorter100|2619_  = \new_Sorter100|2518_  | \new_Sorter100|2519_ ;
  assign \new_Sorter100|2620_  = \new_Sorter100|2520_  & \new_Sorter100|2521_ ;
  assign \new_Sorter100|2621_  = \new_Sorter100|2520_  | \new_Sorter100|2521_ ;
  assign \new_Sorter100|2622_  = \new_Sorter100|2522_  & \new_Sorter100|2523_ ;
  assign \new_Sorter100|2623_  = \new_Sorter100|2522_  | \new_Sorter100|2523_ ;
  assign \new_Sorter100|2624_  = \new_Sorter100|2524_  & \new_Sorter100|2525_ ;
  assign \new_Sorter100|2625_  = \new_Sorter100|2524_  | \new_Sorter100|2525_ ;
  assign \new_Sorter100|2626_  = \new_Sorter100|2526_  & \new_Sorter100|2527_ ;
  assign \new_Sorter100|2627_  = \new_Sorter100|2526_  | \new_Sorter100|2527_ ;
  assign \new_Sorter100|2628_  = \new_Sorter100|2528_  & \new_Sorter100|2529_ ;
  assign \new_Sorter100|2629_  = \new_Sorter100|2528_  | \new_Sorter100|2529_ ;
  assign \new_Sorter100|2630_  = \new_Sorter100|2530_  & \new_Sorter100|2531_ ;
  assign \new_Sorter100|2631_  = \new_Sorter100|2530_  | \new_Sorter100|2531_ ;
  assign \new_Sorter100|2632_  = \new_Sorter100|2532_  & \new_Sorter100|2533_ ;
  assign \new_Sorter100|2633_  = \new_Sorter100|2532_  | \new_Sorter100|2533_ ;
  assign \new_Sorter100|2634_  = \new_Sorter100|2534_  & \new_Sorter100|2535_ ;
  assign \new_Sorter100|2635_  = \new_Sorter100|2534_  | \new_Sorter100|2535_ ;
  assign \new_Sorter100|2636_  = \new_Sorter100|2536_  & \new_Sorter100|2537_ ;
  assign \new_Sorter100|2637_  = \new_Sorter100|2536_  | \new_Sorter100|2537_ ;
  assign \new_Sorter100|2638_  = \new_Sorter100|2538_  & \new_Sorter100|2539_ ;
  assign \new_Sorter100|2639_  = \new_Sorter100|2538_  | \new_Sorter100|2539_ ;
  assign \new_Sorter100|2640_  = \new_Sorter100|2540_  & \new_Sorter100|2541_ ;
  assign \new_Sorter100|2641_  = \new_Sorter100|2540_  | \new_Sorter100|2541_ ;
  assign \new_Sorter100|2642_  = \new_Sorter100|2542_  & \new_Sorter100|2543_ ;
  assign \new_Sorter100|2643_  = \new_Sorter100|2542_  | \new_Sorter100|2543_ ;
  assign \new_Sorter100|2644_  = \new_Sorter100|2544_  & \new_Sorter100|2545_ ;
  assign \new_Sorter100|2645_  = \new_Sorter100|2544_  | \new_Sorter100|2545_ ;
  assign \new_Sorter100|2646_  = \new_Sorter100|2546_  & \new_Sorter100|2547_ ;
  assign \new_Sorter100|2647_  = \new_Sorter100|2546_  | \new_Sorter100|2547_ ;
  assign \new_Sorter100|2648_  = \new_Sorter100|2548_  & \new_Sorter100|2549_ ;
  assign \new_Sorter100|2649_  = \new_Sorter100|2548_  | \new_Sorter100|2549_ ;
  assign \new_Sorter100|2650_  = \new_Sorter100|2550_  & \new_Sorter100|2551_ ;
  assign \new_Sorter100|2651_  = \new_Sorter100|2550_  | \new_Sorter100|2551_ ;
  assign \new_Sorter100|2652_  = \new_Sorter100|2552_  & \new_Sorter100|2553_ ;
  assign \new_Sorter100|2653_  = \new_Sorter100|2552_  | \new_Sorter100|2553_ ;
  assign \new_Sorter100|2654_  = \new_Sorter100|2554_  & \new_Sorter100|2555_ ;
  assign \new_Sorter100|2655_  = \new_Sorter100|2554_  | \new_Sorter100|2555_ ;
  assign \new_Sorter100|2656_  = \new_Sorter100|2556_  & \new_Sorter100|2557_ ;
  assign \new_Sorter100|2657_  = \new_Sorter100|2556_  | \new_Sorter100|2557_ ;
  assign \new_Sorter100|2658_  = \new_Sorter100|2558_  & \new_Sorter100|2559_ ;
  assign \new_Sorter100|2659_  = \new_Sorter100|2558_  | \new_Sorter100|2559_ ;
  assign \new_Sorter100|2660_  = \new_Sorter100|2560_  & \new_Sorter100|2561_ ;
  assign \new_Sorter100|2661_  = \new_Sorter100|2560_  | \new_Sorter100|2561_ ;
  assign \new_Sorter100|2662_  = \new_Sorter100|2562_  & \new_Sorter100|2563_ ;
  assign \new_Sorter100|2663_  = \new_Sorter100|2562_  | \new_Sorter100|2563_ ;
  assign \new_Sorter100|2664_  = \new_Sorter100|2564_  & \new_Sorter100|2565_ ;
  assign \new_Sorter100|2665_  = \new_Sorter100|2564_  | \new_Sorter100|2565_ ;
  assign \new_Sorter100|2666_  = \new_Sorter100|2566_  & \new_Sorter100|2567_ ;
  assign \new_Sorter100|2667_  = \new_Sorter100|2566_  | \new_Sorter100|2567_ ;
  assign \new_Sorter100|2668_  = \new_Sorter100|2568_  & \new_Sorter100|2569_ ;
  assign \new_Sorter100|2669_  = \new_Sorter100|2568_  | \new_Sorter100|2569_ ;
  assign \new_Sorter100|2670_  = \new_Sorter100|2570_  & \new_Sorter100|2571_ ;
  assign \new_Sorter100|2671_  = \new_Sorter100|2570_  | \new_Sorter100|2571_ ;
  assign \new_Sorter100|2672_  = \new_Sorter100|2572_  & \new_Sorter100|2573_ ;
  assign \new_Sorter100|2673_  = \new_Sorter100|2572_  | \new_Sorter100|2573_ ;
  assign \new_Sorter100|2674_  = \new_Sorter100|2574_  & \new_Sorter100|2575_ ;
  assign \new_Sorter100|2675_  = \new_Sorter100|2574_  | \new_Sorter100|2575_ ;
  assign \new_Sorter100|2676_  = \new_Sorter100|2576_  & \new_Sorter100|2577_ ;
  assign \new_Sorter100|2677_  = \new_Sorter100|2576_  | \new_Sorter100|2577_ ;
  assign \new_Sorter100|2678_  = \new_Sorter100|2578_  & \new_Sorter100|2579_ ;
  assign \new_Sorter100|2679_  = \new_Sorter100|2578_  | \new_Sorter100|2579_ ;
  assign \new_Sorter100|2680_  = \new_Sorter100|2580_  & \new_Sorter100|2581_ ;
  assign \new_Sorter100|2681_  = \new_Sorter100|2580_  | \new_Sorter100|2581_ ;
  assign \new_Sorter100|2682_  = \new_Sorter100|2582_  & \new_Sorter100|2583_ ;
  assign \new_Sorter100|2683_  = \new_Sorter100|2582_  | \new_Sorter100|2583_ ;
  assign \new_Sorter100|2684_  = \new_Sorter100|2584_  & \new_Sorter100|2585_ ;
  assign \new_Sorter100|2685_  = \new_Sorter100|2584_  | \new_Sorter100|2585_ ;
  assign \new_Sorter100|2686_  = \new_Sorter100|2586_  & \new_Sorter100|2587_ ;
  assign \new_Sorter100|2687_  = \new_Sorter100|2586_  | \new_Sorter100|2587_ ;
  assign \new_Sorter100|2688_  = \new_Sorter100|2588_  & \new_Sorter100|2589_ ;
  assign \new_Sorter100|2689_  = \new_Sorter100|2588_  | \new_Sorter100|2589_ ;
  assign \new_Sorter100|2690_  = \new_Sorter100|2590_  & \new_Sorter100|2591_ ;
  assign \new_Sorter100|2691_  = \new_Sorter100|2590_  | \new_Sorter100|2591_ ;
  assign \new_Sorter100|2692_  = \new_Sorter100|2592_  & \new_Sorter100|2593_ ;
  assign \new_Sorter100|2693_  = \new_Sorter100|2592_  | \new_Sorter100|2593_ ;
  assign \new_Sorter100|2694_  = \new_Sorter100|2594_  & \new_Sorter100|2595_ ;
  assign \new_Sorter100|2695_  = \new_Sorter100|2594_  | \new_Sorter100|2595_ ;
  assign \new_Sorter100|2696_  = \new_Sorter100|2596_  & \new_Sorter100|2597_ ;
  assign \new_Sorter100|2697_  = \new_Sorter100|2596_  | \new_Sorter100|2597_ ;
  assign \new_Sorter100|2698_  = \new_Sorter100|2598_  & \new_Sorter100|2599_ ;
  assign \new_Sorter100|2699_  = \new_Sorter100|2598_  | \new_Sorter100|2599_ ;
  assign \new_Sorter100|2700_  = \new_Sorter100|2600_ ;
  assign \new_Sorter100|2799_  = \new_Sorter100|2699_ ;
  assign \new_Sorter100|2701_  = \new_Sorter100|2601_  & \new_Sorter100|2602_ ;
  assign \new_Sorter100|2702_  = \new_Sorter100|2601_  | \new_Sorter100|2602_ ;
  assign \new_Sorter100|2703_  = \new_Sorter100|2603_  & \new_Sorter100|2604_ ;
  assign \new_Sorter100|2704_  = \new_Sorter100|2603_  | \new_Sorter100|2604_ ;
  assign \new_Sorter100|2705_  = \new_Sorter100|2605_  & \new_Sorter100|2606_ ;
  assign \new_Sorter100|2706_  = \new_Sorter100|2605_  | \new_Sorter100|2606_ ;
  assign \new_Sorter100|2707_  = \new_Sorter100|2607_  & \new_Sorter100|2608_ ;
  assign \new_Sorter100|2708_  = \new_Sorter100|2607_  | \new_Sorter100|2608_ ;
  assign \new_Sorter100|2709_  = \new_Sorter100|2609_  & \new_Sorter100|2610_ ;
  assign \new_Sorter100|2710_  = \new_Sorter100|2609_  | \new_Sorter100|2610_ ;
  assign \new_Sorter100|2711_  = \new_Sorter100|2611_  & \new_Sorter100|2612_ ;
  assign \new_Sorter100|2712_  = \new_Sorter100|2611_  | \new_Sorter100|2612_ ;
  assign \new_Sorter100|2713_  = \new_Sorter100|2613_  & \new_Sorter100|2614_ ;
  assign \new_Sorter100|2714_  = \new_Sorter100|2613_  | \new_Sorter100|2614_ ;
  assign \new_Sorter100|2715_  = \new_Sorter100|2615_  & \new_Sorter100|2616_ ;
  assign \new_Sorter100|2716_  = \new_Sorter100|2615_  | \new_Sorter100|2616_ ;
  assign \new_Sorter100|2717_  = \new_Sorter100|2617_  & \new_Sorter100|2618_ ;
  assign \new_Sorter100|2718_  = \new_Sorter100|2617_  | \new_Sorter100|2618_ ;
  assign \new_Sorter100|2719_  = \new_Sorter100|2619_  & \new_Sorter100|2620_ ;
  assign \new_Sorter100|2720_  = \new_Sorter100|2619_  | \new_Sorter100|2620_ ;
  assign \new_Sorter100|2721_  = \new_Sorter100|2621_  & \new_Sorter100|2622_ ;
  assign \new_Sorter100|2722_  = \new_Sorter100|2621_  | \new_Sorter100|2622_ ;
  assign \new_Sorter100|2723_  = \new_Sorter100|2623_  & \new_Sorter100|2624_ ;
  assign \new_Sorter100|2724_  = \new_Sorter100|2623_  | \new_Sorter100|2624_ ;
  assign \new_Sorter100|2725_  = \new_Sorter100|2625_  & \new_Sorter100|2626_ ;
  assign \new_Sorter100|2726_  = \new_Sorter100|2625_  | \new_Sorter100|2626_ ;
  assign \new_Sorter100|2727_  = \new_Sorter100|2627_  & \new_Sorter100|2628_ ;
  assign \new_Sorter100|2728_  = \new_Sorter100|2627_  | \new_Sorter100|2628_ ;
  assign \new_Sorter100|2729_  = \new_Sorter100|2629_  & \new_Sorter100|2630_ ;
  assign \new_Sorter100|2730_  = \new_Sorter100|2629_  | \new_Sorter100|2630_ ;
  assign \new_Sorter100|2731_  = \new_Sorter100|2631_  & \new_Sorter100|2632_ ;
  assign \new_Sorter100|2732_  = \new_Sorter100|2631_  | \new_Sorter100|2632_ ;
  assign \new_Sorter100|2733_  = \new_Sorter100|2633_  & \new_Sorter100|2634_ ;
  assign \new_Sorter100|2734_  = \new_Sorter100|2633_  | \new_Sorter100|2634_ ;
  assign \new_Sorter100|2735_  = \new_Sorter100|2635_  & \new_Sorter100|2636_ ;
  assign \new_Sorter100|2736_  = \new_Sorter100|2635_  | \new_Sorter100|2636_ ;
  assign \new_Sorter100|2737_  = \new_Sorter100|2637_  & \new_Sorter100|2638_ ;
  assign \new_Sorter100|2738_  = \new_Sorter100|2637_  | \new_Sorter100|2638_ ;
  assign \new_Sorter100|2739_  = \new_Sorter100|2639_  & \new_Sorter100|2640_ ;
  assign \new_Sorter100|2740_  = \new_Sorter100|2639_  | \new_Sorter100|2640_ ;
  assign \new_Sorter100|2741_  = \new_Sorter100|2641_  & \new_Sorter100|2642_ ;
  assign \new_Sorter100|2742_  = \new_Sorter100|2641_  | \new_Sorter100|2642_ ;
  assign \new_Sorter100|2743_  = \new_Sorter100|2643_  & \new_Sorter100|2644_ ;
  assign \new_Sorter100|2744_  = \new_Sorter100|2643_  | \new_Sorter100|2644_ ;
  assign \new_Sorter100|2745_  = \new_Sorter100|2645_  & \new_Sorter100|2646_ ;
  assign \new_Sorter100|2746_  = \new_Sorter100|2645_  | \new_Sorter100|2646_ ;
  assign \new_Sorter100|2747_  = \new_Sorter100|2647_  & \new_Sorter100|2648_ ;
  assign \new_Sorter100|2748_  = \new_Sorter100|2647_  | \new_Sorter100|2648_ ;
  assign \new_Sorter100|2749_  = \new_Sorter100|2649_  & \new_Sorter100|2650_ ;
  assign \new_Sorter100|2750_  = \new_Sorter100|2649_  | \new_Sorter100|2650_ ;
  assign \new_Sorter100|2751_  = \new_Sorter100|2651_  & \new_Sorter100|2652_ ;
  assign \new_Sorter100|2752_  = \new_Sorter100|2651_  | \new_Sorter100|2652_ ;
  assign \new_Sorter100|2753_  = \new_Sorter100|2653_  & \new_Sorter100|2654_ ;
  assign \new_Sorter100|2754_  = \new_Sorter100|2653_  | \new_Sorter100|2654_ ;
  assign \new_Sorter100|2755_  = \new_Sorter100|2655_  & \new_Sorter100|2656_ ;
  assign \new_Sorter100|2756_  = \new_Sorter100|2655_  | \new_Sorter100|2656_ ;
  assign \new_Sorter100|2757_  = \new_Sorter100|2657_  & \new_Sorter100|2658_ ;
  assign \new_Sorter100|2758_  = \new_Sorter100|2657_  | \new_Sorter100|2658_ ;
  assign \new_Sorter100|2759_  = \new_Sorter100|2659_  & \new_Sorter100|2660_ ;
  assign \new_Sorter100|2760_  = \new_Sorter100|2659_  | \new_Sorter100|2660_ ;
  assign \new_Sorter100|2761_  = \new_Sorter100|2661_  & \new_Sorter100|2662_ ;
  assign \new_Sorter100|2762_  = \new_Sorter100|2661_  | \new_Sorter100|2662_ ;
  assign \new_Sorter100|2763_  = \new_Sorter100|2663_  & \new_Sorter100|2664_ ;
  assign \new_Sorter100|2764_  = \new_Sorter100|2663_  | \new_Sorter100|2664_ ;
  assign \new_Sorter100|2765_  = \new_Sorter100|2665_  & \new_Sorter100|2666_ ;
  assign \new_Sorter100|2766_  = \new_Sorter100|2665_  | \new_Sorter100|2666_ ;
  assign \new_Sorter100|2767_  = \new_Sorter100|2667_  & \new_Sorter100|2668_ ;
  assign \new_Sorter100|2768_  = \new_Sorter100|2667_  | \new_Sorter100|2668_ ;
  assign \new_Sorter100|2769_  = \new_Sorter100|2669_  & \new_Sorter100|2670_ ;
  assign \new_Sorter100|2770_  = \new_Sorter100|2669_  | \new_Sorter100|2670_ ;
  assign \new_Sorter100|2771_  = \new_Sorter100|2671_  & \new_Sorter100|2672_ ;
  assign \new_Sorter100|2772_  = \new_Sorter100|2671_  | \new_Sorter100|2672_ ;
  assign \new_Sorter100|2773_  = \new_Sorter100|2673_  & \new_Sorter100|2674_ ;
  assign \new_Sorter100|2774_  = \new_Sorter100|2673_  | \new_Sorter100|2674_ ;
  assign \new_Sorter100|2775_  = \new_Sorter100|2675_  & \new_Sorter100|2676_ ;
  assign \new_Sorter100|2776_  = \new_Sorter100|2675_  | \new_Sorter100|2676_ ;
  assign \new_Sorter100|2777_  = \new_Sorter100|2677_  & \new_Sorter100|2678_ ;
  assign \new_Sorter100|2778_  = \new_Sorter100|2677_  | \new_Sorter100|2678_ ;
  assign \new_Sorter100|2779_  = \new_Sorter100|2679_  & \new_Sorter100|2680_ ;
  assign \new_Sorter100|2780_  = \new_Sorter100|2679_  | \new_Sorter100|2680_ ;
  assign \new_Sorter100|2781_  = \new_Sorter100|2681_  & \new_Sorter100|2682_ ;
  assign \new_Sorter100|2782_  = \new_Sorter100|2681_  | \new_Sorter100|2682_ ;
  assign \new_Sorter100|2783_  = \new_Sorter100|2683_  & \new_Sorter100|2684_ ;
  assign \new_Sorter100|2784_  = \new_Sorter100|2683_  | \new_Sorter100|2684_ ;
  assign \new_Sorter100|2785_  = \new_Sorter100|2685_  & \new_Sorter100|2686_ ;
  assign \new_Sorter100|2786_  = \new_Sorter100|2685_  | \new_Sorter100|2686_ ;
  assign \new_Sorter100|2787_  = \new_Sorter100|2687_  & \new_Sorter100|2688_ ;
  assign \new_Sorter100|2788_  = \new_Sorter100|2687_  | \new_Sorter100|2688_ ;
  assign \new_Sorter100|2789_  = \new_Sorter100|2689_  & \new_Sorter100|2690_ ;
  assign \new_Sorter100|2790_  = \new_Sorter100|2689_  | \new_Sorter100|2690_ ;
  assign \new_Sorter100|2791_  = \new_Sorter100|2691_  & \new_Sorter100|2692_ ;
  assign \new_Sorter100|2792_  = \new_Sorter100|2691_  | \new_Sorter100|2692_ ;
  assign \new_Sorter100|2793_  = \new_Sorter100|2693_  & \new_Sorter100|2694_ ;
  assign \new_Sorter100|2794_  = \new_Sorter100|2693_  | \new_Sorter100|2694_ ;
  assign \new_Sorter100|2795_  = \new_Sorter100|2695_  & \new_Sorter100|2696_ ;
  assign \new_Sorter100|2796_  = \new_Sorter100|2695_  | \new_Sorter100|2696_ ;
  assign \new_Sorter100|2797_  = \new_Sorter100|2697_  & \new_Sorter100|2698_ ;
  assign \new_Sorter100|2798_  = \new_Sorter100|2697_  | \new_Sorter100|2698_ ;
  assign \new_Sorter100|2800_  = \new_Sorter100|2700_  & \new_Sorter100|2701_ ;
  assign \new_Sorter100|2801_  = \new_Sorter100|2700_  | \new_Sorter100|2701_ ;
  assign \new_Sorter100|2802_  = \new_Sorter100|2702_  & \new_Sorter100|2703_ ;
  assign \new_Sorter100|2803_  = \new_Sorter100|2702_  | \new_Sorter100|2703_ ;
  assign \new_Sorter100|2804_  = \new_Sorter100|2704_  & \new_Sorter100|2705_ ;
  assign \new_Sorter100|2805_  = \new_Sorter100|2704_  | \new_Sorter100|2705_ ;
  assign \new_Sorter100|2806_  = \new_Sorter100|2706_  & \new_Sorter100|2707_ ;
  assign \new_Sorter100|2807_  = \new_Sorter100|2706_  | \new_Sorter100|2707_ ;
  assign \new_Sorter100|2808_  = \new_Sorter100|2708_  & \new_Sorter100|2709_ ;
  assign \new_Sorter100|2809_  = \new_Sorter100|2708_  | \new_Sorter100|2709_ ;
  assign \new_Sorter100|2810_  = \new_Sorter100|2710_  & \new_Sorter100|2711_ ;
  assign \new_Sorter100|2811_  = \new_Sorter100|2710_  | \new_Sorter100|2711_ ;
  assign \new_Sorter100|2812_  = \new_Sorter100|2712_  & \new_Sorter100|2713_ ;
  assign \new_Sorter100|2813_  = \new_Sorter100|2712_  | \new_Sorter100|2713_ ;
  assign \new_Sorter100|2814_  = \new_Sorter100|2714_  & \new_Sorter100|2715_ ;
  assign \new_Sorter100|2815_  = \new_Sorter100|2714_  | \new_Sorter100|2715_ ;
  assign \new_Sorter100|2816_  = \new_Sorter100|2716_  & \new_Sorter100|2717_ ;
  assign \new_Sorter100|2817_  = \new_Sorter100|2716_  | \new_Sorter100|2717_ ;
  assign \new_Sorter100|2818_  = \new_Sorter100|2718_  & \new_Sorter100|2719_ ;
  assign \new_Sorter100|2819_  = \new_Sorter100|2718_  | \new_Sorter100|2719_ ;
  assign \new_Sorter100|2820_  = \new_Sorter100|2720_  & \new_Sorter100|2721_ ;
  assign \new_Sorter100|2821_  = \new_Sorter100|2720_  | \new_Sorter100|2721_ ;
  assign \new_Sorter100|2822_  = \new_Sorter100|2722_  & \new_Sorter100|2723_ ;
  assign \new_Sorter100|2823_  = \new_Sorter100|2722_  | \new_Sorter100|2723_ ;
  assign \new_Sorter100|2824_  = \new_Sorter100|2724_  & \new_Sorter100|2725_ ;
  assign \new_Sorter100|2825_  = \new_Sorter100|2724_  | \new_Sorter100|2725_ ;
  assign \new_Sorter100|2826_  = \new_Sorter100|2726_  & \new_Sorter100|2727_ ;
  assign \new_Sorter100|2827_  = \new_Sorter100|2726_  | \new_Sorter100|2727_ ;
  assign \new_Sorter100|2828_  = \new_Sorter100|2728_  & \new_Sorter100|2729_ ;
  assign \new_Sorter100|2829_  = \new_Sorter100|2728_  | \new_Sorter100|2729_ ;
  assign \new_Sorter100|2830_  = \new_Sorter100|2730_  & \new_Sorter100|2731_ ;
  assign \new_Sorter100|2831_  = \new_Sorter100|2730_  | \new_Sorter100|2731_ ;
  assign \new_Sorter100|2832_  = \new_Sorter100|2732_  & \new_Sorter100|2733_ ;
  assign \new_Sorter100|2833_  = \new_Sorter100|2732_  | \new_Sorter100|2733_ ;
  assign \new_Sorter100|2834_  = \new_Sorter100|2734_  & \new_Sorter100|2735_ ;
  assign \new_Sorter100|2835_  = \new_Sorter100|2734_  | \new_Sorter100|2735_ ;
  assign \new_Sorter100|2836_  = \new_Sorter100|2736_  & \new_Sorter100|2737_ ;
  assign \new_Sorter100|2837_  = \new_Sorter100|2736_  | \new_Sorter100|2737_ ;
  assign \new_Sorter100|2838_  = \new_Sorter100|2738_  & \new_Sorter100|2739_ ;
  assign \new_Sorter100|2839_  = \new_Sorter100|2738_  | \new_Sorter100|2739_ ;
  assign \new_Sorter100|2840_  = \new_Sorter100|2740_  & \new_Sorter100|2741_ ;
  assign \new_Sorter100|2841_  = \new_Sorter100|2740_  | \new_Sorter100|2741_ ;
  assign \new_Sorter100|2842_  = \new_Sorter100|2742_  & \new_Sorter100|2743_ ;
  assign \new_Sorter100|2843_  = \new_Sorter100|2742_  | \new_Sorter100|2743_ ;
  assign \new_Sorter100|2844_  = \new_Sorter100|2744_  & \new_Sorter100|2745_ ;
  assign \new_Sorter100|2845_  = \new_Sorter100|2744_  | \new_Sorter100|2745_ ;
  assign \new_Sorter100|2846_  = \new_Sorter100|2746_  & \new_Sorter100|2747_ ;
  assign \new_Sorter100|2847_  = \new_Sorter100|2746_  | \new_Sorter100|2747_ ;
  assign \new_Sorter100|2848_  = \new_Sorter100|2748_  & \new_Sorter100|2749_ ;
  assign \new_Sorter100|2849_  = \new_Sorter100|2748_  | \new_Sorter100|2749_ ;
  assign \new_Sorter100|2850_  = \new_Sorter100|2750_  & \new_Sorter100|2751_ ;
  assign \new_Sorter100|2851_  = \new_Sorter100|2750_  | \new_Sorter100|2751_ ;
  assign \new_Sorter100|2852_  = \new_Sorter100|2752_  & \new_Sorter100|2753_ ;
  assign \new_Sorter100|2853_  = \new_Sorter100|2752_  | \new_Sorter100|2753_ ;
  assign \new_Sorter100|2854_  = \new_Sorter100|2754_  & \new_Sorter100|2755_ ;
  assign \new_Sorter100|2855_  = \new_Sorter100|2754_  | \new_Sorter100|2755_ ;
  assign \new_Sorter100|2856_  = \new_Sorter100|2756_  & \new_Sorter100|2757_ ;
  assign \new_Sorter100|2857_  = \new_Sorter100|2756_  | \new_Sorter100|2757_ ;
  assign \new_Sorter100|2858_  = \new_Sorter100|2758_  & \new_Sorter100|2759_ ;
  assign \new_Sorter100|2859_  = \new_Sorter100|2758_  | \new_Sorter100|2759_ ;
  assign \new_Sorter100|2860_  = \new_Sorter100|2760_  & \new_Sorter100|2761_ ;
  assign \new_Sorter100|2861_  = \new_Sorter100|2760_  | \new_Sorter100|2761_ ;
  assign \new_Sorter100|2862_  = \new_Sorter100|2762_  & \new_Sorter100|2763_ ;
  assign \new_Sorter100|2863_  = \new_Sorter100|2762_  | \new_Sorter100|2763_ ;
  assign \new_Sorter100|2864_  = \new_Sorter100|2764_  & \new_Sorter100|2765_ ;
  assign \new_Sorter100|2865_  = \new_Sorter100|2764_  | \new_Sorter100|2765_ ;
  assign \new_Sorter100|2866_  = \new_Sorter100|2766_  & \new_Sorter100|2767_ ;
  assign \new_Sorter100|2867_  = \new_Sorter100|2766_  | \new_Sorter100|2767_ ;
  assign \new_Sorter100|2868_  = \new_Sorter100|2768_  & \new_Sorter100|2769_ ;
  assign \new_Sorter100|2869_  = \new_Sorter100|2768_  | \new_Sorter100|2769_ ;
  assign \new_Sorter100|2870_  = \new_Sorter100|2770_  & \new_Sorter100|2771_ ;
  assign \new_Sorter100|2871_  = \new_Sorter100|2770_  | \new_Sorter100|2771_ ;
  assign \new_Sorter100|2872_  = \new_Sorter100|2772_  & \new_Sorter100|2773_ ;
  assign \new_Sorter100|2873_  = \new_Sorter100|2772_  | \new_Sorter100|2773_ ;
  assign \new_Sorter100|2874_  = \new_Sorter100|2774_  & \new_Sorter100|2775_ ;
  assign \new_Sorter100|2875_  = \new_Sorter100|2774_  | \new_Sorter100|2775_ ;
  assign \new_Sorter100|2876_  = \new_Sorter100|2776_  & \new_Sorter100|2777_ ;
  assign \new_Sorter100|2877_  = \new_Sorter100|2776_  | \new_Sorter100|2777_ ;
  assign \new_Sorter100|2878_  = \new_Sorter100|2778_  & \new_Sorter100|2779_ ;
  assign \new_Sorter100|2879_  = \new_Sorter100|2778_  | \new_Sorter100|2779_ ;
  assign \new_Sorter100|2880_  = \new_Sorter100|2780_  & \new_Sorter100|2781_ ;
  assign \new_Sorter100|2881_  = \new_Sorter100|2780_  | \new_Sorter100|2781_ ;
  assign \new_Sorter100|2882_  = \new_Sorter100|2782_  & \new_Sorter100|2783_ ;
  assign \new_Sorter100|2883_  = \new_Sorter100|2782_  | \new_Sorter100|2783_ ;
  assign \new_Sorter100|2884_  = \new_Sorter100|2784_  & \new_Sorter100|2785_ ;
  assign \new_Sorter100|2885_  = \new_Sorter100|2784_  | \new_Sorter100|2785_ ;
  assign \new_Sorter100|2886_  = \new_Sorter100|2786_  & \new_Sorter100|2787_ ;
  assign \new_Sorter100|2887_  = \new_Sorter100|2786_  | \new_Sorter100|2787_ ;
  assign \new_Sorter100|2888_  = \new_Sorter100|2788_  & \new_Sorter100|2789_ ;
  assign \new_Sorter100|2889_  = \new_Sorter100|2788_  | \new_Sorter100|2789_ ;
  assign \new_Sorter100|2890_  = \new_Sorter100|2790_  & \new_Sorter100|2791_ ;
  assign \new_Sorter100|2891_  = \new_Sorter100|2790_  | \new_Sorter100|2791_ ;
  assign \new_Sorter100|2892_  = \new_Sorter100|2792_  & \new_Sorter100|2793_ ;
  assign \new_Sorter100|2893_  = \new_Sorter100|2792_  | \new_Sorter100|2793_ ;
  assign \new_Sorter100|2894_  = \new_Sorter100|2794_  & \new_Sorter100|2795_ ;
  assign \new_Sorter100|2895_  = \new_Sorter100|2794_  | \new_Sorter100|2795_ ;
  assign \new_Sorter100|2896_  = \new_Sorter100|2796_  & \new_Sorter100|2797_ ;
  assign \new_Sorter100|2897_  = \new_Sorter100|2796_  | \new_Sorter100|2797_ ;
  assign \new_Sorter100|2898_  = \new_Sorter100|2798_  & \new_Sorter100|2799_ ;
  assign \new_Sorter100|2899_  = \new_Sorter100|2798_  | \new_Sorter100|2799_ ;
  assign \new_Sorter100|2900_  = \new_Sorter100|2800_ ;
  assign \new_Sorter100|2999_  = \new_Sorter100|2899_ ;
  assign \new_Sorter100|2901_  = \new_Sorter100|2801_  & \new_Sorter100|2802_ ;
  assign \new_Sorter100|2902_  = \new_Sorter100|2801_  | \new_Sorter100|2802_ ;
  assign \new_Sorter100|2903_  = \new_Sorter100|2803_  & \new_Sorter100|2804_ ;
  assign \new_Sorter100|2904_  = \new_Sorter100|2803_  | \new_Sorter100|2804_ ;
  assign \new_Sorter100|2905_  = \new_Sorter100|2805_  & \new_Sorter100|2806_ ;
  assign \new_Sorter100|2906_  = \new_Sorter100|2805_  | \new_Sorter100|2806_ ;
  assign \new_Sorter100|2907_  = \new_Sorter100|2807_  & \new_Sorter100|2808_ ;
  assign \new_Sorter100|2908_  = \new_Sorter100|2807_  | \new_Sorter100|2808_ ;
  assign \new_Sorter100|2909_  = \new_Sorter100|2809_  & \new_Sorter100|2810_ ;
  assign \new_Sorter100|2910_  = \new_Sorter100|2809_  | \new_Sorter100|2810_ ;
  assign \new_Sorter100|2911_  = \new_Sorter100|2811_  & \new_Sorter100|2812_ ;
  assign \new_Sorter100|2912_  = \new_Sorter100|2811_  | \new_Sorter100|2812_ ;
  assign \new_Sorter100|2913_  = \new_Sorter100|2813_  & \new_Sorter100|2814_ ;
  assign \new_Sorter100|2914_  = \new_Sorter100|2813_  | \new_Sorter100|2814_ ;
  assign \new_Sorter100|2915_  = \new_Sorter100|2815_  & \new_Sorter100|2816_ ;
  assign \new_Sorter100|2916_  = \new_Sorter100|2815_  | \new_Sorter100|2816_ ;
  assign \new_Sorter100|2917_  = \new_Sorter100|2817_  & \new_Sorter100|2818_ ;
  assign \new_Sorter100|2918_  = \new_Sorter100|2817_  | \new_Sorter100|2818_ ;
  assign \new_Sorter100|2919_  = \new_Sorter100|2819_  & \new_Sorter100|2820_ ;
  assign \new_Sorter100|2920_  = \new_Sorter100|2819_  | \new_Sorter100|2820_ ;
  assign \new_Sorter100|2921_  = \new_Sorter100|2821_  & \new_Sorter100|2822_ ;
  assign \new_Sorter100|2922_  = \new_Sorter100|2821_  | \new_Sorter100|2822_ ;
  assign \new_Sorter100|2923_  = \new_Sorter100|2823_  & \new_Sorter100|2824_ ;
  assign \new_Sorter100|2924_  = \new_Sorter100|2823_  | \new_Sorter100|2824_ ;
  assign \new_Sorter100|2925_  = \new_Sorter100|2825_  & \new_Sorter100|2826_ ;
  assign \new_Sorter100|2926_  = \new_Sorter100|2825_  | \new_Sorter100|2826_ ;
  assign \new_Sorter100|2927_  = \new_Sorter100|2827_  & \new_Sorter100|2828_ ;
  assign \new_Sorter100|2928_  = \new_Sorter100|2827_  | \new_Sorter100|2828_ ;
  assign \new_Sorter100|2929_  = \new_Sorter100|2829_  & \new_Sorter100|2830_ ;
  assign \new_Sorter100|2930_  = \new_Sorter100|2829_  | \new_Sorter100|2830_ ;
  assign \new_Sorter100|2931_  = \new_Sorter100|2831_  & \new_Sorter100|2832_ ;
  assign \new_Sorter100|2932_  = \new_Sorter100|2831_  | \new_Sorter100|2832_ ;
  assign \new_Sorter100|2933_  = \new_Sorter100|2833_  & \new_Sorter100|2834_ ;
  assign \new_Sorter100|2934_  = \new_Sorter100|2833_  | \new_Sorter100|2834_ ;
  assign \new_Sorter100|2935_  = \new_Sorter100|2835_  & \new_Sorter100|2836_ ;
  assign \new_Sorter100|2936_  = \new_Sorter100|2835_  | \new_Sorter100|2836_ ;
  assign \new_Sorter100|2937_  = \new_Sorter100|2837_  & \new_Sorter100|2838_ ;
  assign \new_Sorter100|2938_  = \new_Sorter100|2837_  | \new_Sorter100|2838_ ;
  assign \new_Sorter100|2939_  = \new_Sorter100|2839_  & \new_Sorter100|2840_ ;
  assign \new_Sorter100|2940_  = \new_Sorter100|2839_  | \new_Sorter100|2840_ ;
  assign \new_Sorter100|2941_  = \new_Sorter100|2841_  & \new_Sorter100|2842_ ;
  assign \new_Sorter100|2942_  = \new_Sorter100|2841_  | \new_Sorter100|2842_ ;
  assign \new_Sorter100|2943_  = \new_Sorter100|2843_  & \new_Sorter100|2844_ ;
  assign \new_Sorter100|2944_  = \new_Sorter100|2843_  | \new_Sorter100|2844_ ;
  assign \new_Sorter100|2945_  = \new_Sorter100|2845_  & \new_Sorter100|2846_ ;
  assign \new_Sorter100|2946_  = \new_Sorter100|2845_  | \new_Sorter100|2846_ ;
  assign \new_Sorter100|2947_  = \new_Sorter100|2847_  & \new_Sorter100|2848_ ;
  assign \new_Sorter100|2948_  = \new_Sorter100|2847_  | \new_Sorter100|2848_ ;
  assign \new_Sorter100|2949_  = \new_Sorter100|2849_  & \new_Sorter100|2850_ ;
  assign \new_Sorter100|2950_  = \new_Sorter100|2849_  | \new_Sorter100|2850_ ;
  assign \new_Sorter100|2951_  = \new_Sorter100|2851_  & \new_Sorter100|2852_ ;
  assign \new_Sorter100|2952_  = \new_Sorter100|2851_  | \new_Sorter100|2852_ ;
  assign \new_Sorter100|2953_  = \new_Sorter100|2853_  & \new_Sorter100|2854_ ;
  assign \new_Sorter100|2954_  = \new_Sorter100|2853_  | \new_Sorter100|2854_ ;
  assign \new_Sorter100|2955_  = \new_Sorter100|2855_  & \new_Sorter100|2856_ ;
  assign \new_Sorter100|2956_  = \new_Sorter100|2855_  | \new_Sorter100|2856_ ;
  assign \new_Sorter100|2957_  = \new_Sorter100|2857_  & \new_Sorter100|2858_ ;
  assign \new_Sorter100|2958_  = \new_Sorter100|2857_  | \new_Sorter100|2858_ ;
  assign \new_Sorter100|2959_  = \new_Sorter100|2859_  & \new_Sorter100|2860_ ;
  assign \new_Sorter100|2960_  = \new_Sorter100|2859_  | \new_Sorter100|2860_ ;
  assign \new_Sorter100|2961_  = \new_Sorter100|2861_  & \new_Sorter100|2862_ ;
  assign \new_Sorter100|2962_  = \new_Sorter100|2861_  | \new_Sorter100|2862_ ;
  assign \new_Sorter100|2963_  = \new_Sorter100|2863_  & \new_Sorter100|2864_ ;
  assign \new_Sorter100|2964_  = \new_Sorter100|2863_  | \new_Sorter100|2864_ ;
  assign \new_Sorter100|2965_  = \new_Sorter100|2865_  & \new_Sorter100|2866_ ;
  assign \new_Sorter100|2966_  = \new_Sorter100|2865_  | \new_Sorter100|2866_ ;
  assign \new_Sorter100|2967_  = \new_Sorter100|2867_  & \new_Sorter100|2868_ ;
  assign \new_Sorter100|2968_  = \new_Sorter100|2867_  | \new_Sorter100|2868_ ;
  assign \new_Sorter100|2969_  = \new_Sorter100|2869_  & \new_Sorter100|2870_ ;
  assign \new_Sorter100|2970_  = \new_Sorter100|2869_  | \new_Sorter100|2870_ ;
  assign \new_Sorter100|2971_  = \new_Sorter100|2871_  & \new_Sorter100|2872_ ;
  assign \new_Sorter100|2972_  = \new_Sorter100|2871_  | \new_Sorter100|2872_ ;
  assign \new_Sorter100|2973_  = \new_Sorter100|2873_  & \new_Sorter100|2874_ ;
  assign \new_Sorter100|2974_  = \new_Sorter100|2873_  | \new_Sorter100|2874_ ;
  assign \new_Sorter100|2975_  = \new_Sorter100|2875_  & \new_Sorter100|2876_ ;
  assign \new_Sorter100|2976_  = \new_Sorter100|2875_  | \new_Sorter100|2876_ ;
  assign \new_Sorter100|2977_  = \new_Sorter100|2877_  & \new_Sorter100|2878_ ;
  assign \new_Sorter100|2978_  = \new_Sorter100|2877_  | \new_Sorter100|2878_ ;
  assign \new_Sorter100|2979_  = \new_Sorter100|2879_  & \new_Sorter100|2880_ ;
  assign \new_Sorter100|2980_  = \new_Sorter100|2879_  | \new_Sorter100|2880_ ;
  assign \new_Sorter100|2981_  = \new_Sorter100|2881_  & \new_Sorter100|2882_ ;
  assign \new_Sorter100|2982_  = \new_Sorter100|2881_  | \new_Sorter100|2882_ ;
  assign \new_Sorter100|2983_  = \new_Sorter100|2883_  & \new_Sorter100|2884_ ;
  assign \new_Sorter100|2984_  = \new_Sorter100|2883_  | \new_Sorter100|2884_ ;
  assign \new_Sorter100|2985_  = \new_Sorter100|2885_  & \new_Sorter100|2886_ ;
  assign \new_Sorter100|2986_  = \new_Sorter100|2885_  | \new_Sorter100|2886_ ;
  assign \new_Sorter100|2987_  = \new_Sorter100|2887_  & \new_Sorter100|2888_ ;
  assign \new_Sorter100|2988_  = \new_Sorter100|2887_  | \new_Sorter100|2888_ ;
  assign \new_Sorter100|2989_  = \new_Sorter100|2889_  & \new_Sorter100|2890_ ;
  assign \new_Sorter100|2990_  = \new_Sorter100|2889_  | \new_Sorter100|2890_ ;
  assign \new_Sorter100|2991_  = \new_Sorter100|2891_  & \new_Sorter100|2892_ ;
  assign \new_Sorter100|2992_  = \new_Sorter100|2891_  | \new_Sorter100|2892_ ;
  assign \new_Sorter100|2993_  = \new_Sorter100|2893_  & \new_Sorter100|2894_ ;
  assign \new_Sorter100|2994_  = \new_Sorter100|2893_  | \new_Sorter100|2894_ ;
  assign \new_Sorter100|2995_  = \new_Sorter100|2895_  & \new_Sorter100|2896_ ;
  assign \new_Sorter100|2996_  = \new_Sorter100|2895_  | \new_Sorter100|2896_ ;
  assign \new_Sorter100|2997_  = \new_Sorter100|2897_  & \new_Sorter100|2898_ ;
  assign \new_Sorter100|2998_  = \new_Sorter100|2897_  | \new_Sorter100|2898_ ;
  assign \new_Sorter100|3000_  = \new_Sorter100|2900_  & \new_Sorter100|2901_ ;
  assign \new_Sorter100|3001_  = \new_Sorter100|2900_  | \new_Sorter100|2901_ ;
  assign \new_Sorter100|3002_  = \new_Sorter100|2902_  & \new_Sorter100|2903_ ;
  assign \new_Sorter100|3003_  = \new_Sorter100|2902_  | \new_Sorter100|2903_ ;
  assign \new_Sorter100|3004_  = \new_Sorter100|2904_  & \new_Sorter100|2905_ ;
  assign \new_Sorter100|3005_  = \new_Sorter100|2904_  | \new_Sorter100|2905_ ;
  assign \new_Sorter100|3006_  = \new_Sorter100|2906_  & \new_Sorter100|2907_ ;
  assign \new_Sorter100|3007_  = \new_Sorter100|2906_  | \new_Sorter100|2907_ ;
  assign \new_Sorter100|3008_  = \new_Sorter100|2908_  & \new_Sorter100|2909_ ;
  assign \new_Sorter100|3009_  = \new_Sorter100|2908_  | \new_Sorter100|2909_ ;
  assign \new_Sorter100|3010_  = \new_Sorter100|2910_  & \new_Sorter100|2911_ ;
  assign \new_Sorter100|3011_  = \new_Sorter100|2910_  | \new_Sorter100|2911_ ;
  assign \new_Sorter100|3012_  = \new_Sorter100|2912_  & \new_Sorter100|2913_ ;
  assign \new_Sorter100|3013_  = \new_Sorter100|2912_  | \new_Sorter100|2913_ ;
  assign \new_Sorter100|3014_  = \new_Sorter100|2914_  & \new_Sorter100|2915_ ;
  assign \new_Sorter100|3015_  = \new_Sorter100|2914_  | \new_Sorter100|2915_ ;
  assign \new_Sorter100|3016_  = \new_Sorter100|2916_  & \new_Sorter100|2917_ ;
  assign \new_Sorter100|3017_  = \new_Sorter100|2916_  | \new_Sorter100|2917_ ;
  assign \new_Sorter100|3018_  = \new_Sorter100|2918_  & \new_Sorter100|2919_ ;
  assign \new_Sorter100|3019_  = \new_Sorter100|2918_  | \new_Sorter100|2919_ ;
  assign \new_Sorter100|3020_  = \new_Sorter100|2920_  & \new_Sorter100|2921_ ;
  assign \new_Sorter100|3021_  = \new_Sorter100|2920_  | \new_Sorter100|2921_ ;
  assign \new_Sorter100|3022_  = \new_Sorter100|2922_  & \new_Sorter100|2923_ ;
  assign \new_Sorter100|3023_  = \new_Sorter100|2922_  | \new_Sorter100|2923_ ;
  assign \new_Sorter100|3024_  = \new_Sorter100|2924_  & \new_Sorter100|2925_ ;
  assign \new_Sorter100|3025_  = \new_Sorter100|2924_  | \new_Sorter100|2925_ ;
  assign \new_Sorter100|3026_  = \new_Sorter100|2926_  & \new_Sorter100|2927_ ;
  assign \new_Sorter100|3027_  = \new_Sorter100|2926_  | \new_Sorter100|2927_ ;
  assign \new_Sorter100|3028_  = \new_Sorter100|2928_  & \new_Sorter100|2929_ ;
  assign \new_Sorter100|3029_  = \new_Sorter100|2928_  | \new_Sorter100|2929_ ;
  assign \new_Sorter100|3030_  = \new_Sorter100|2930_  & \new_Sorter100|2931_ ;
  assign \new_Sorter100|3031_  = \new_Sorter100|2930_  | \new_Sorter100|2931_ ;
  assign \new_Sorter100|3032_  = \new_Sorter100|2932_  & \new_Sorter100|2933_ ;
  assign \new_Sorter100|3033_  = \new_Sorter100|2932_  | \new_Sorter100|2933_ ;
  assign \new_Sorter100|3034_  = \new_Sorter100|2934_  & \new_Sorter100|2935_ ;
  assign \new_Sorter100|3035_  = \new_Sorter100|2934_  | \new_Sorter100|2935_ ;
  assign \new_Sorter100|3036_  = \new_Sorter100|2936_  & \new_Sorter100|2937_ ;
  assign \new_Sorter100|3037_  = \new_Sorter100|2936_  | \new_Sorter100|2937_ ;
  assign \new_Sorter100|3038_  = \new_Sorter100|2938_  & \new_Sorter100|2939_ ;
  assign \new_Sorter100|3039_  = \new_Sorter100|2938_  | \new_Sorter100|2939_ ;
  assign \new_Sorter100|3040_  = \new_Sorter100|2940_  & \new_Sorter100|2941_ ;
  assign \new_Sorter100|3041_  = \new_Sorter100|2940_  | \new_Sorter100|2941_ ;
  assign \new_Sorter100|3042_  = \new_Sorter100|2942_  & \new_Sorter100|2943_ ;
  assign \new_Sorter100|3043_  = \new_Sorter100|2942_  | \new_Sorter100|2943_ ;
  assign \new_Sorter100|3044_  = \new_Sorter100|2944_  & \new_Sorter100|2945_ ;
  assign \new_Sorter100|3045_  = \new_Sorter100|2944_  | \new_Sorter100|2945_ ;
  assign \new_Sorter100|3046_  = \new_Sorter100|2946_  & \new_Sorter100|2947_ ;
  assign \new_Sorter100|3047_  = \new_Sorter100|2946_  | \new_Sorter100|2947_ ;
  assign \new_Sorter100|3048_  = \new_Sorter100|2948_  & \new_Sorter100|2949_ ;
  assign \new_Sorter100|3049_  = \new_Sorter100|2948_  | \new_Sorter100|2949_ ;
  assign \new_Sorter100|3050_  = \new_Sorter100|2950_  & \new_Sorter100|2951_ ;
  assign \new_Sorter100|3051_  = \new_Sorter100|2950_  | \new_Sorter100|2951_ ;
  assign \new_Sorter100|3052_  = \new_Sorter100|2952_  & \new_Sorter100|2953_ ;
  assign \new_Sorter100|3053_  = \new_Sorter100|2952_  | \new_Sorter100|2953_ ;
  assign \new_Sorter100|3054_  = \new_Sorter100|2954_  & \new_Sorter100|2955_ ;
  assign \new_Sorter100|3055_  = \new_Sorter100|2954_  | \new_Sorter100|2955_ ;
  assign \new_Sorter100|3056_  = \new_Sorter100|2956_  & \new_Sorter100|2957_ ;
  assign \new_Sorter100|3057_  = \new_Sorter100|2956_  | \new_Sorter100|2957_ ;
  assign \new_Sorter100|3058_  = \new_Sorter100|2958_  & \new_Sorter100|2959_ ;
  assign \new_Sorter100|3059_  = \new_Sorter100|2958_  | \new_Sorter100|2959_ ;
  assign \new_Sorter100|3060_  = \new_Sorter100|2960_  & \new_Sorter100|2961_ ;
  assign \new_Sorter100|3061_  = \new_Sorter100|2960_  | \new_Sorter100|2961_ ;
  assign \new_Sorter100|3062_  = \new_Sorter100|2962_  & \new_Sorter100|2963_ ;
  assign \new_Sorter100|3063_  = \new_Sorter100|2962_  | \new_Sorter100|2963_ ;
  assign \new_Sorter100|3064_  = \new_Sorter100|2964_  & \new_Sorter100|2965_ ;
  assign \new_Sorter100|3065_  = \new_Sorter100|2964_  | \new_Sorter100|2965_ ;
  assign \new_Sorter100|3066_  = \new_Sorter100|2966_  & \new_Sorter100|2967_ ;
  assign \new_Sorter100|3067_  = \new_Sorter100|2966_  | \new_Sorter100|2967_ ;
  assign \new_Sorter100|3068_  = \new_Sorter100|2968_  & \new_Sorter100|2969_ ;
  assign \new_Sorter100|3069_  = \new_Sorter100|2968_  | \new_Sorter100|2969_ ;
  assign \new_Sorter100|3070_  = \new_Sorter100|2970_  & \new_Sorter100|2971_ ;
  assign \new_Sorter100|3071_  = \new_Sorter100|2970_  | \new_Sorter100|2971_ ;
  assign \new_Sorter100|3072_  = \new_Sorter100|2972_  & \new_Sorter100|2973_ ;
  assign \new_Sorter100|3073_  = \new_Sorter100|2972_  | \new_Sorter100|2973_ ;
  assign \new_Sorter100|3074_  = \new_Sorter100|2974_  & \new_Sorter100|2975_ ;
  assign \new_Sorter100|3075_  = \new_Sorter100|2974_  | \new_Sorter100|2975_ ;
  assign \new_Sorter100|3076_  = \new_Sorter100|2976_  & \new_Sorter100|2977_ ;
  assign \new_Sorter100|3077_  = \new_Sorter100|2976_  | \new_Sorter100|2977_ ;
  assign \new_Sorter100|3078_  = \new_Sorter100|2978_  & \new_Sorter100|2979_ ;
  assign \new_Sorter100|3079_  = \new_Sorter100|2978_  | \new_Sorter100|2979_ ;
  assign \new_Sorter100|3080_  = \new_Sorter100|2980_  & \new_Sorter100|2981_ ;
  assign \new_Sorter100|3081_  = \new_Sorter100|2980_  | \new_Sorter100|2981_ ;
  assign \new_Sorter100|3082_  = \new_Sorter100|2982_  & \new_Sorter100|2983_ ;
  assign \new_Sorter100|3083_  = \new_Sorter100|2982_  | \new_Sorter100|2983_ ;
  assign \new_Sorter100|3084_  = \new_Sorter100|2984_  & \new_Sorter100|2985_ ;
  assign \new_Sorter100|3085_  = \new_Sorter100|2984_  | \new_Sorter100|2985_ ;
  assign \new_Sorter100|3086_  = \new_Sorter100|2986_  & \new_Sorter100|2987_ ;
  assign \new_Sorter100|3087_  = \new_Sorter100|2986_  | \new_Sorter100|2987_ ;
  assign \new_Sorter100|3088_  = \new_Sorter100|2988_  & \new_Sorter100|2989_ ;
  assign \new_Sorter100|3089_  = \new_Sorter100|2988_  | \new_Sorter100|2989_ ;
  assign \new_Sorter100|3090_  = \new_Sorter100|2990_  & \new_Sorter100|2991_ ;
  assign \new_Sorter100|3091_  = \new_Sorter100|2990_  | \new_Sorter100|2991_ ;
  assign \new_Sorter100|3092_  = \new_Sorter100|2992_  & \new_Sorter100|2993_ ;
  assign \new_Sorter100|3093_  = \new_Sorter100|2992_  | \new_Sorter100|2993_ ;
  assign \new_Sorter100|3094_  = \new_Sorter100|2994_  & \new_Sorter100|2995_ ;
  assign \new_Sorter100|3095_  = \new_Sorter100|2994_  | \new_Sorter100|2995_ ;
  assign \new_Sorter100|3096_  = \new_Sorter100|2996_  & \new_Sorter100|2997_ ;
  assign \new_Sorter100|3097_  = \new_Sorter100|2996_  | \new_Sorter100|2997_ ;
  assign \new_Sorter100|3098_  = \new_Sorter100|2998_  & \new_Sorter100|2999_ ;
  assign \new_Sorter100|3099_  = \new_Sorter100|2998_  | \new_Sorter100|2999_ ;
  assign \new_Sorter100|3100_  = \new_Sorter100|3000_ ;
  assign \new_Sorter100|3199_  = \new_Sorter100|3099_ ;
  assign \new_Sorter100|3101_  = \new_Sorter100|3001_  & \new_Sorter100|3002_ ;
  assign \new_Sorter100|3102_  = \new_Sorter100|3001_  | \new_Sorter100|3002_ ;
  assign \new_Sorter100|3103_  = \new_Sorter100|3003_  & \new_Sorter100|3004_ ;
  assign \new_Sorter100|3104_  = \new_Sorter100|3003_  | \new_Sorter100|3004_ ;
  assign \new_Sorter100|3105_  = \new_Sorter100|3005_  & \new_Sorter100|3006_ ;
  assign \new_Sorter100|3106_  = \new_Sorter100|3005_  | \new_Sorter100|3006_ ;
  assign \new_Sorter100|3107_  = \new_Sorter100|3007_  & \new_Sorter100|3008_ ;
  assign \new_Sorter100|3108_  = \new_Sorter100|3007_  | \new_Sorter100|3008_ ;
  assign \new_Sorter100|3109_  = \new_Sorter100|3009_  & \new_Sorter100|3010_ ;
  assign \new_Sorter100|3110_  = \new_Sorter100|3009_  | \new_Sorter100|3010_ ;
  assign \new_Sorter100|3111_  = \new_Sorter100|3011_  & \new_Sorter100|3012_ ;
  assign \new_Sorter100|3112_  = \new_Sorter100|3011_  | \new_Sorter100|3012_ ;
  assign \new_Sorter100|3113_  = \new_Sorter100|3013_  & \new_Sorter100|3014_ ;
  assign \new_Sorter100|3114_  = \new_Sorter100|3013_  | \new_Sorter100|3014_ ;
  assign \new_Sorter100|3115_  = \new_Sorter100|3015_  & \new_Sorter100|3016_ ;
  assign \new_Sorter100|3116_  = \new_Sorter100|3015_  | \new_Sorter100|3016_ ;
  assign \new_Sorter100|3117_  = \new_Sorter100|3017_  & \new_Sorter100|3018_ ;
  assign \new_Sorter100|3118_  = \new_Sorter100|3017_  | \new_Sorter100|3018_ ;
  assign \new_Sorter100|3119_  = \new_Sorter100|3019_  & \new_Sorter100|3020_ ;
  assign \new_Sorter100|3120_  = \new_Sorter100|3019_  | \new_Sorter100|3020_ ;
  assign \new_Sorter100|3121_  = \new_Sorter100|3021_  & \new_Sorter100|3022_ ;
  assign \new_Sorter100|3122_  = \new_Sorter100|3021_  | \new_Sorter100|3022_ ;
  assign \new_Sorter100|3123_  = \new_Sorter100|3023_  & \new_Sorter100|3024_ ;
  assign \new_Sorter100|3124_  = \new_Sorter100|3023_  | \new_Sorter100|3024_ ;
  assign \new_Sorter100|3125_  = \new_Sorter100|3025_  & \new_Sorter100|3026_ ;
  assign \new_Sorter100|3126_  = \new_Sorter100|3025_  | \new_Sorter100|3026_ ;
  assign \new_Sorter100|3127_  = \new_Sorter100|3027_  & \new_Sorter100|3028_ ;
  assign \new_Sorter100|3128_  = \new_Sorter100|3027_  | \new_Sorter100|3028_ ;
  assign \new_Sorter100|3129_  = \new_Sorter100|3029_  & \new_Sorter100|3030_ ;
  assign \new_Sorter100|3130_  = \new_Sorter100|3029_  | \new_Sorter100|3030_ ;
  assign \new_Sorter100|3131_  = \new_Sorter100|3031_  & \new_Sorter100|3032_ ;
  assign \new_Sorter100|3132_  = \new_Sorter100|3031_  | \new_Sorter100|3032_ ;
  assign \new_Sorter100|3133_  = \new_Sorter100|3033_  & \new_Sorter100|3034_ ;
  assign \new_Sorter100|3134_  = \new_Sorter100|3033_  | \new_Sorter100|3034_ ;
  assign \new_Sorter100|3135_  = \new_Sorter100|3035_  & \new_Sorter100|3036_ ;
  assign \new_Sorter100|3136_  = \new_Sorter100|3035_  | \new_Sorter100|3036_ ;
  assign \new_Sorter100|3137_  = \new_Sorter100|3037_  & \new_Sorter100|3038_ ;
  assign \new_Sorter100|3138_  = \new_Sorter100|3037_  | \new_Sorter100|3038_ ;
  assign \new_Sorter100|3139_  = \new_Sorter100|3039_  & \new_Sorter100|3040_ ;
  assign \new_Sorter100|3140_  = \new_Sorter100|3039_  | \new_Sorter100|3040_ ;
  assign \new_Sorter100|3141_  = \new_Sorter100|3041_  & \new_Sorter100|3042_ ;
  assign \new_Sorter100|3142_  = \new_Sorter100|3041_  | \new_Sorter100|3042_ ;
  assign \new_Sorter100|3143_  = \new_Sorter100|3043_  & \new_Sorter100|3044_ ;
  assign \new_Sorter100|3144_  = \new_Sorter100|3043_  | \new_Sorter100|3044_ ;
  assign \new_Sorter100|3145_  = \new_Sorter100|3045_  & \new_Sorter100|3046_ ;
  assign \new_Sorter100|3146_  = \new_Sorter100|3045_  | \new_Sorter100|3046_ ;
  assign \new_Sorter100|3147_  = \new_Sorter100|3047_  & \new_Sorter100|3048_ ;
  assign \new_Sorter100|3148_  = \new_Sorter100|3047_  | \new_Sorter100|3048_ ;
  assign \new_Sorter100|3149_  = \new_Sorter100|3049_  & \new_Sorter100|3050_ ;
  assign \new_Sorter100|3150_  = \new_Sorter100|3049_  | \new_Sorter100|3050_ ;
  assign \new_Sorter100|3151_  = \new_Sorter100|3051_  & \new_Sorter100|3052_ ;
  assign \new_Sorter100|3152_  = \new_Sorter100|3051_  | \new_Sorter100|3052_ ;
  assign \new_Sorter100|3153_  = \new_Sorter100|3053_  & \new_Sorter100|3054_ ;
  assign \new_Sorter100|3154_  = \new_Sorter100|3053_  | \new_Sorter100|3054_ ;
  assign \new_Sorter100|3155_  = \new_Sorter100|3055_  & \new_Sorter100|3056_ ;
  assign \new_Sorter100|3156_  = \new_Sorter100|3055_  | \new_Sorter100|3056_ ;
  assign \new_Sorter100|3157_  = \new_Sorter100|3057_  & \new_Sorter100|3058_ ;
  assign \new_Sorter100|3158_  = \new_Sorter100|3057_  | \new_Sorter100|3058_ ;
  assign \new_Sorter100|3159_  = \new_Sorter100|3059_  & \new_Sorter100|3060_ ;
  assign \new_Sorter100|3160_  = \new_Sorter100|3059_  | \new_Sorter100|3060_ ;
  assign \new_Sorter100|3161_  = \new_Sorter100|3061_  & \new_Sorter100|3062_ ;
  assign \new_Sorter100|3162_  = \new_Sorter100|3061_  | \new_Sorter100|3062_ ;
  assign \new_Sorter100|3163_  = \new_Sorter100|3063_  & \new_Sorter100|3064_ ;
  assign \new_Sorter100|3164_  = \new_Sorter100|3063_  | \new_Sorter100|3064_ ;
  assign \new_Sorter100|3165_  = \new_Sorter100|3065_  & \new_Sorter100|3066_ ;
  assign \new_Sorter100|3166_  = \new_Sorter100|3065_  | \new_Sorter100|3066_ ;
  assign \new_Sorter100|3167_  = \new_Sorter100|3067_  & \new_Sorter100|3068_ ;
  assign \new_Sorter100|3168_  = \new_Sorter100|3067_  | \new_Sorter100|3068_ ;
  assign \new_Sorter100|3169_  = \new_Sorter100|3069_  & \new_Sorter100|3070_ ;
  assign \new_Sorter100|3170_  = \new_Sorter100|3069_  | \new_Sorter100|3070_ ;
  assign \new_Sorter100|3171_  = \new_Sorter100|3071_  & \new_Sorter100|3072_ ;
  assign \new_Sorter100|3172_  = \new_Sorter100|3071_  | \new_Sorter100|3072_ ;
  assign \new_Sorter100|3173_  = \new_Sorter100|3073_  & \new_Sorter100|3074_ ;
  assign \new_Sorter100|3174_  = \new_Sorter100|3073_  | \new_Sorter100|3074_ ;
  assign \new_Sorter100|3175_  = \new_Sorter100|3075_  & \new_Sorter100|3076_ ;
  assign \new_Sorter100|3176_  = \new_Sorter100|3075_  | \new_Sorter100|3076_ ;
  assign \new_Sorter100|3177_  = \new_Sorter100|3077_  & \new_Sorter100|3078_ ;
  assign \new_Sorter100|3178_  = \new_Sorter100|3077_  | \new_Sorter100|3078_ ;
  assign \new_Sorter100|3179_  = \new_Sorter100|3079_  & \new_Sorter100|3080_ ;
  assign \new_Sorter100|3180_  = \new_Sorter100|3079_  | \new_Sorter100|3080_ ;
  assign \new_Sorter100|3181_  = \new_Sorter100|3081_  & \new_Sorter100|3082_ ;
  assign \new_Sorter100|3182_  = \new_Sorter100|3081_  | \new_Sorter100|3082_ ;
  assign \new_Sorter100|3183_  = \new_Sorter100|3083_  & \new_Sorter100|3084_ ;
  assign \new_Sorter100|3184_  = \new_Sorter100|3083_  | \new_Sorter100|3084_ ;
  assign \new_Sorter100|3185_  = \new_Sorter100|3085_  & \new_Sorter100|3086_ ;
  assign \new_Sorter100|3186_  = \new_Sorter100|3085_  | \new_Sorter100|3086_ ;
  assign \new_Sorter100|3187_  = \new_Sorter100|3087_  & \new_Sorter100|3088_ ;
  assign \new_Sorter100|3188_  = \new_Sorter100|3087_  | \new_Sorter100|3088_ ;
  assign \new_Sorter100|3189_  = \new_Sorter100|3089_  & \new_Sorter100|3090_ ;
  assign \new_Sorter100|3190_  = \new_Sorter100|3089_  | \new_Sorter100|3090_ ;
  assign \new_Sorter100|3191_  = \new_Sorter100|3091_  & \new_Sorter100|3092_ ;
  assign \new_Sorter100|3192_  = \new_Sorter100|3091_  | \new_Sorter100|3092_ ;
  assign \new_Sorter100|3193_  = \new_Sorter100|3093_  & \new_Sorter100|3094_ ;
  assign \new_Sorter100|3194_  = \new_Sorter100|3093_  | \new_Sorter100|3094_ ;
  assign \new_Sorter100|3195_  = \new_Sorter100|3095_  & \new_Sorter100|3096_ ;
  assign \new_Sorter100|3196_  = \new_Sorter100|3095_  | \new_Sorter100|3096_ ;
  assign \new_Sorter100|3197_  = \new_Sorter100|3097_  & \new_Sorter100|3098_ ;
  assign \new_Sorter100|3198_  = \new_Sorter100|3097_  | \new_Sorter100|3098_ ;
  assign \new_Sorter100|3200_  = \new_Sorter100|3100_  & \new_Sorter100|3101_ ;
  assign \new_Sorter100|3201_  = \new_Sorter100|3100_  | \new_Sorter100|3101_ ;
  assign \new_Sorter100|3202_  = \new_Sorter100|3102_  & \new_Sorter100|3103_ ;
  assign \new_Sorter100|3203_  = \new_Sorter100|3102_  | \new_Sorter100|3103_ ;
  assign \new_Sorter100|3204_  = \new_Sorter100|3104_  & \new_Sorter100|3105_ ;
  assign \new_Sorter100|3205_  = \new_Sorter100|3104_  | \new_Sorter100|3105_ ;
  assign \new_Sorter100|3206_  = \new_Sorter100|3106_  & \new_Sorter100|3107_ ;
  assign \new_Sorter100|3207_  = \new_Sorter100|3106_  | \new_Sorter100|3107_ ;
  assign \new_Sorter100|3208_  = \new_Sorter100|3108_  & \new_Sorter100|3109_ ;
  assign \new_Sorter100|3209_  = \new_Sorter100|3108_  | \new_Sorter100|3109_ ;
  assign \new_Sorter100|3210_  = \new_Sorter100|3110_  & \new_Sorter100|3111_ ;
  assign \new_Sorter100|3211_  = \new_Sorter100|3110_  | \new_Sorter100|3111_ ;
  assign \new_Sorter100|3212_  = \new_Sorter100|3112_  & \new_Sorter100|3113_ ;
  assign \new_Sorter100|3213_  = \new_Sorter100|3112_  | \new_Sorter100|3113_ ;
  assign \new_Sorter100|3214_  = \new_Sorter100|3114_  & \new_Sorter100|3115_ ;
  assign \new_Sorter100|3215_  = \new_Sorter100|3114_  | \new_Sorter100|3115_ ;
  assign \new_Sorter100|3216_  = \new_Sorter100|3116_  & \new_Sorter100|3117_ ;
  assign \new_Sorter100|3217_  = \new_Sorter100|3116_  | \new_Sorter100|3117_ ;
  assign \new_Sorter100|3218_  = \new_Sorter100|3118_  & \new_Sorter100|3119_ ;
  assign \new_Sorter100|3219_  = \new_Sorter100|3118_  | \new_Sorter100|3119_ ;
  assign \new_Sorter100|3220_  = \new_Sorter100|3120_  & \new_Sorter100|3121_ ;
  assign \new_Sorter100|3221_  = \new_Sorter100|3120_  | \new_Sorter100|3121_ ;
  assign \new_Sorter100|3222_  = \new_Sorter100|3122_  & \new_Sorter100|3123_ ;
  assign \new_Sorter100|3223_  = \new_Sorter100|3122_  | \new_Sorter100|3123_ ;
  assign \new_Sorter100|3224_  = \new_Sorter100|3124_  & \new_Sorter100|3125_ ;
  assign \new_Sorter100|3225_  = \new_Sorter100|3124_  | \new_Sorter100|3125_ ;
  assign \new_Sorter100|3226_  = \new_Sorter100|3126_  & \new_Sorter100|3127_ ;
  assign \new_Sorter100|3227_  = \new_Sorter100|3126_  | \new_Sorter100|3127_ ;
  assign \new_Sorter100|3228_  = \new_Sorter100|3128_  & \new_Sorter100|3129_ ;
  assign \new_Sorter100|3229_  = \new_Sorter100|3128_  | \new_Sorter100|3129_ ;
  assign \new_Sorter100|3230_  = \new_Sorter100|3130_  & \new_Sorter100|3131_ ;
  assign \new_Sorter100|3231_  = \new_Sorter100|3130_  | \new_Sorter100|3131_ ;
  assign \new_Sorter100|3232_  = \new_Sorter100|3132_  & \new_Sorter100|3133_ ;
  assign \new_Sorter100|3233_  = \new_Sorter100|3132_  | \new_Sorter100|3133_ ;
  assign \new_Sorter100|3234_  = \new_Sorter100|3134_  & \new_Sorter100|3135_ ;
  assign \new_Sorter100|3235_  = \new_Sorter100|3134_  | \new_Sorter100|3135_ ;
  assign \new_Sorter100|3236_  = \new_Sorter100|3136_  & \new_Sorter100|3137_ ;
  assign \new_Sorter100|3237_  = \new_Sorter100|3136_  | \new_Sorter100|3137_ ;
  assign \new_Sorter100|3238_  = \new_Sorter100|3138_  & \new_Sorter100|3139_ ;
  assign \new_Sorter100|3239_  = \new_Sorter100|3138_  | \new_Sorter100|3139_ ;
  assign \new_Sorter100|3240_  = \new_Sorter100|3140_  & \new_Sorter100|3141_ ;
  assign \new_Sorter100|3241_  = \new_Sorter100|3140_  | \new_Sorter100|3141_ ;
  assign \new_Sorter100|3242_  = \new_Sorter100|3142_  & \new_Sorter100|3143_ ;
  assign \new_Sorter100|3243_  = \new_Sorter100|3142_  | \new_Sorter100|3143_ ;
  assign \new_Sorter100|3244_  = \new_Sorter100|3144_  & \new_Sorter100|3145_ ;
  assign \new_Sorter100|3245_  = \new_Sorter100|3144_  | \new_Sorter100|3145_ ;
  assign \new_Sorter100|3246_  = \new_Sorter100|3146_  & \new_Sorter100|3147_ ;
  assign \new_Sorter100|3247_  = \new_Sorter100|3146_  | \new_Sorter100|3147_ ;
  assign \new_Sorter100|3248_  = \new_Sorter100|3148_  & \new_Sorter100|3149_ ;
  assign \new_Sorter100|3249_  = \new_Sorter100|3148_  | \new_Sorter100|3149_ ;
  assign \new_Sorter100|3250_  = \new_Sorter100|3150_  & \new_Sorter100|3151_ ;
  assign \new_Sorter100|3251_  = \new_Sorter100|3150_  | \new_Sorter100|3151_ ;
  assign \new_Sorter100|3252_  = \new_Sorter100|3152_  & \new_Sorter100|3153_ ;
  assign \new_Sorter100|3253_  = \new_Sorter100|3152_  | \new_Sorter100|3153_ ;
  assign \new_Sorter100|3254_  = \new_Sorter100|3154_  & \new_Sorter100|3155_ ;
  assign \new_Sorter100|3255_  = \new_Sorter100|3154_  | \new_Sorter100|3155_ ;
  assign \new_Sorter100|3256_  = \new_Sorter100|3156_  & \new_Sorter100|3157_ ;
  assign \new_Sorter100|3257_  = \new_Sorter100|3156_  | \new_Sorter100|3157_ ;
  assign \new_Sorter100|3258_  = \new_Sorter100|3158_  & \new_Sorter100|3159_ ;
  assign \new_Sorter100|3259_  = \new_Sorter100|3158_  | \new_Sorter100|3159_ ;
  assign \new_Sorter100|3260_  = \new_Sorter100|3160_  & \new_Sorter100|3161_ ;
  assign \new_Sorter100|3261_  = \new_Sorter100|3160_  | \new_Sorter100|3161_ ;
  assign \new_Sorter100|3262_  = \new_Sorter100|3162_  & \new_Sorter100|3163_ ;
  assign \new_Sorter100|3263_  = \new_Sorter100|3162_  | \new_Sorter100|3163_ ;
  assign \new_Sorter100|3264_  = \new_Sorter100|3164_  & \new_Sorter100|3165_ ;
  assign \new_Sorter100|3265_  = \new_Sorter100|3164_  | \new_Sorter100|3165_ ;
  assign \new_Sorter100|3266_  = \new_Sorter100|3166_  & \new_Sorter100|3167_ ;
  assign \new_Sorter100|3267_  = \new_Sorter100|3166_  | \new_Sorter100|3167_ ;
  assign \new_Sorter100|3268_  = \new_Sorter100|3168_  & \new_Sorter100|3169_ ;
  assign \new_Sorter100|3269_  = \new_Sorter100|3168_  | \new_Sorter100|3169_ ;
  assign \new_Sorter100|3270_  = \new_Sorter100|3170_  & \new_Sorter100|3171_ ;
  assign \new_Sorter100|3271_  = \new_Sorter100|3170_  | \new_Sorter100|3171_ ;
  assign \new_Sorter100|3272_  = \new_Sorter100|3172_  & \new_Sorter100|3173_ ;
  assign \new_Sorter100|3273_  = \new_Sorter100|3172_  | \new_Sorter100|3173_ ;
  assign \new_Sorter100|3274_  = \new_Sorter100|3174_  & \new_Sorter100|3175_ ;
  assign \new_Sorter100|3275_  = \new_Sorter100|3174_  | \new_Sorter100|3175_ ;
  assign \new_Sorter100|3276_  = \new_Sorter100|3176_  & \new_Sorter100|3177_ ;
  assign \new_Sorter100|3277_  = \new_Sorter100|3176_  | \new_Sorter100|3177_ ;
  assign \new_Sorter100|3278_  = \new_Sorter100|3178_  & \new_Sorter100|3179_ ;
  assign \new_Sorter100|3279_  = \new_Sorter100|3178_  | \new_Sorter100|3179_ ;
  assign \new_Sorter100|3280_  = \new_Sorter100|3180_  & \new_Sorter100|3181_ ;
  assign \new_Sorter100|3281_  = \new_Sorter100|3180_  | \new_Sorter100|3181_ ;
  assign \new_Sorter100|3282_  = \new_Sorter100|3182_  & \new_Sorter100|3183_ ;
  assign \new_Sorter100|3283_  = \new_Sorter100|3182_  | \new_Sorter100|3183_ ;
  assign \new_Sorter100|3284_  = \new_Sorter100|3184_  & \new_Sorter100|3185_ ;
  assign \new_Sorter100|3285_  = \new_Sorter100|3184_  | \new_Sorter100|3185_ ;
  assign \new_Sorter100|3286_  = \new_Sorter100|3186_  & \new_Sorter100|3187_ ;
  assign \new_Sorter100|3287_  = \new_Sorter100|3186_  | \new_Sorter100|3187_ ;
  assign \new_Sorter100|3288_  = \new_Sorter100|3188_  & \new_Sorter100|3189_ ;
  assign \new_Sorter100|3289_  = \new_Sorter100|3188_  | \new_Sorter100|3189_ ;
  assign \new_Sorter100|3290_  = \new_Sorter100|3190_  & \new_Sorter100|3191_ ;
  assign \new_Sorter100|3291_  = \new_Sorter100|3190_  | \new_Sorter100|3191_ ;
  assign \new_Sorter100|3292_  = \new_Sorter100|3192_  & \new_Sorter100|3193_ ;
  assign \new_Sorter100|3293_  = \new_Sorter100|3192_  | \new_Sorter100|3193_ ;
  assign \new_Sorter100|3294_  = \new_Sorter100|3194_  & \new_Sorter100|3195_ ;
  assign \new_Sorter100|3295_  = \new_Sorter100|3194_  | \new_Sorter100|3195_ ;
  assign \new_Sorter100|3296_  = \new_Sorter100|3196_  & \new_Sorter100|3197_ ;
  assign \new_Sorter100|3297_  = \new_Sorter100|3196_  | \new_Sorter100|3197_ ;
  assign \new_Sorter100|3298_  = \new_Sorter100|3198_  & \new_Sorter100|3199_ ;
  assign \new_Sorter100|3299_  = \new_Sorter100|3198_  | \new_Sorter100|3199_ ;
  assign \new_Sorter100|3300_  = \new_Sorter100|3200_ ;
  assign \new_Sorter100|3399_  = \new_Sorter100|3299_ ;
  assign \new_Sorter100|3301_  = \new_Sorter100|3201_  & \new_Sorter100|3202_ ;
  assign \new_Sorter100|3302_  = \new_Sorter100|3201_  | \new_Sorter100|3202_ ;
  assign \new_Sorter100|3303_  = \new_Sorter100|3203_  & \new_Sorter100|3204_ ;
  assign \new_Sorter100|3304_  = \new_Sorter100|3203_  | \new_Sorter100|3204_ ;
  assign \new_Sorter100|3305_  = \new_Sorter100|3205_  & \new_Sorter100|3206_ ;
  assign \new_Sorter100|3306_  = \new_Sorter100|3205_  | \new_Sorter100|3206_ ;
  assign \new_Sorter100|3307_  = \new_Sorter100|3207_  & \new_Sorter100|3208_ ;
  assign \new_Sorter100|3308_  = \new_Sorter100|3207_  | \new_Sorter100|3208_ ;
  assign \new_Sorter100|3309_  = \new_Sorter100|3209_  & \new_Sorter100|3210_ ;
  assign \new_Sorter100|3310_  = \new_Sorter100|3209_  | \new_Sorter100|3210_ ;
  assign \new_Sorter100|3311_  = \new_Sorter100|3211_  & \new_Sorter100|3212_ ;
  assign \new_Sorter100|3312_  = \new_Sorter100|3211_  | \new_Sorter100|3212_ ;
  assign \new_Sorter100|3313_  = \new_Sorter100|3213_  & \new_Sorter100|3214_ ;
  assign \new_Sorter100|3314_  = \new_Sorter100|3213_  | \new_Sorter100|3214_ ;
  assign \new_Sorter100|3315_  = \new_Sorter100|3215_  & \new_Sorter100|3216_ ;
  assign \new_Sorter100|3316_  = \new_Sorter100|3215_  | \new_Sorter100|3216_ ;
  assign \new_Sorter100|3317_  = \new_Sorter100|3217_  & \new_Sorter100|3218_ ;
  assign \new_Sorter100|3318_  = \new_Sorter100|3217_  | \new_Sorter100|3218_ ;
  assign \new_Sorter100|3319_  = \new_Sorter100|3219_  & \new_Sorter100|3220_ ;
  assign \new_Sorter100|3320_  = \new_Sorter100|3219_  | \new_Sorter100|3220_ ;
  assign \new_Sorter100|3321_  = \new_Sorter100|3221_  & \new_Sorter100|3222_ ;
  assign \new_Sorter100|3322_  = \new_Sorter100|3221_  | \new_Sorter100|3222_ ;
  assign \new_Sorter100|3323_  = \new_Sorter100|3223_  & \new_Sorter100|3224_ ;
  assign \new_Sorter100|3324_  = \new_Sorter100|3223_  | \new_Sorter100|3224_ ;
  assign \new_Sorter100|3325_  = \new_Sorter100|3225_  & \new_Sorter100|3226_ ;
  assign \new_Sorter100|3326_  = \new_Sorter100|3225_  | \new_Sorter100|3226_ ;
  assign \new_Sorter100|3327_  = \new_Sorter100|3227_  & \new_Sorter100|3228_ ;
  assign \new_Sorter100|3328_  = \new_Sorter100|3227_  | \new_Sorter100|3228_ ;
  assign \new_Sorter100|3329_  = \new_Sorter100|3229_  & \new_Sorter100|3230_ ;
  assign \new_Sorter100|3330_  = \new_Sorter100|3229_  | \new_Sorter100|3230_ ;
  assign \new_Sorter100|3331_  = \new_Sorter100|3231_  & \new_Sorter100|3232_ ;
  assign \new_Sorter100|3332_  = \new_Sorter100|3231_  | \new_Sorter100|3232_ ;
  assign \new_Sorter100|3333_  = \new_Sorter100|3233_  & \new_Sorter100|3234_ ;
  assign \new_Sorter100|3334_  = \new_Sorter100|3233_  | \new_Sorter100|3234_ ;
  assign \new_Sorter100|3335_  = \new_Sorter100|3235_  & \new_Sorter100|3236_ ;
  assign \new_Sorter100|3336_  = \new_Sorter100|3235_  | \new_Sorter100|3236_ ;
  assign \new_Sorter100|3337_  = \new_Sorter100|3237_  & \new_Sorter100|3238_ ;
  assign \new_Sorter100|3338_  = \new_Sorter100|3237_  | \new_Sorter100|3238_ ;
  assign \new_Sorter100|3339_  = \new_Sorter100|3239_  & \new_Sorter100|3240_ ;
  assign \new_Sorter100|3340_  = \new_Sorter100|3239_  | \new_Sorter100|3240_ ;
  assign \new_Sorter100|3341_  = \new_Sorter100|3241_  & \new_Sorter100|3242_ ;
  assign \new_Sorter100|3342_  = \new_Sorter100|3241_  | \new_Sorter100|3242_ ;
  assign \new_Sorter100|3343_  = \new_Sorter100|3243_  & \new_Sorter100|3244_ ;
  assign \new_Sorter100|3344_  = \new_Sorter100|3243_  | \new_Sorter100|3244_ ;
  assign \new_Sorter100|3345_  = \new_Sorter100|3245_  & \new_Sorter100|3246_ ;
  assign \new_Sorter100|3346_  = \new_Sorter100|3245_  | \new_Sorter100|3246_ ;
  assign \new_Sorter100|3347_  = \new_Sorter100|3247_  & \new_Sorter100|3248_ ;
  assign \new_Sorter100|3348_  = \new_Sorter100|3247_  | \new_Sorter100|3248_ ;
  assign \new_Sorter100|3349_  = \new_Sorter100|3249_  & \new_Sorter100|3250_ ;
  assign \new_Sorter100|3350_  = \new_Sorter100|3249_  | \new_Sorter100|3250_ ;
  assign \new_Sorter100|3351_  = \new_Sorter100|3251_  & \new_Sorter100|3252_ ;
  assign \new_Sorter100|3352_  = \new_Sorter100|3251_  | \new_Sorter100|3252_ ;
  assign \new_Sorter100|3353_  = \new_Sorter100|3253_  & \new_Sorter100|3254_ ;
  assign \new_Sorter100|3354_  = \new_Sorter100|3253_  | \new_Sorter100|3254_ ;
  assign \new_Sorter100|3355_  = \new_Sorter100|3255_  & \new_Sorter100|3256_ ;
  assign \new_Sorter100|3356_  = \new_Sorter100|3255_  | \new_Sorter100|3256_ ;
  assign \new_Sorter100|3357_  = \new_Sorter100|3257_  & \new_Sorter100|3258_ ;
  assign \new_Sorter100|3358_  = \new_Sorter100|3257_  | \new_Sorter100|3258_ ;
  assign \new_Sorter100|3359_  = \new_Sorter100|3259_  & \new_Sorter100|3260_ ;
  assign \new_Sorter100|3360_  = \new_Sorter100|3259_  | \new_Sorter100|3260_ ;
  assign \new_Sorter100|3361_  = \new_Sorter100|3261_  & \new_Sorter100|3262_ ;
  assign \new_Sorter100|3362_  = \new_Sorter100|3261_  | \new_Sorter100|3262_ ;
  assign \new_Sorter100|3363_  = \new_Sorter100|3263_  & \new_Sorter100|3264_ ;
  assign \new_Sorter100|3364_  = \new_Sorter100|3263_  | \new_Sorter100|3264_ ;
  assign \new_Sorter100|3365_  = \new_Sorter100|3265_  & \new_Sorter100|3266_ ;
  assign \new_Sorter100|3366_  = \new_Sorter100|3265_  | \new_Sorter100|3266_ ;
  assign \new_Sorter100|3367_  = \new_Sorter100|3267_  & \new_Sorter100|3268_ ;
  assign \new_Sorter100|3368_  = \new_Sorter100|3267_  | \new_Sorter100|3268_ ;
  assign \new_Sorter100|3369_  = \new_Sorter100|3269_  & \new_Sorter100|3270_ ;
  assign \new_Sorter100|3370_  = \new_Sorter100|3269_  | \new_Sorter100|3270_ ;
  assign \new_Sorter100|3371_  = \new_Sorter100|3271_  & \new_Sorter100|3272_ ;
  assign \new_Sorter100|3372_  = \new_Sorter100|3271_  | \new_Sorter100|3272_ ;
  assign \new_Sorter100|3373_  = \new_Sorter100|3273_  & \new_Sorter100|3274_ ;
  assign \new_Sorter100|3374_  = \new_Sorter100|3273_  | \new_Sorter100|3274_ ;
  assign \new_Sorter100|3375_  = \new_Sorter100|3275_  & \new_Sorter100|3276_ ;
  assign \new_Sorter100|3376_  = \new_Sorter100|3275_  | \new_Sorter100|3276_ ;
  assign \new_Sorter100|3377_  = \new_Sorter100|3277_  & \new_Sorter100|3278_ ;
  assign \new_Sorter100|3378_  = \new_Sorter100|3277_  | \new_Sorter100|3278_ ;
  assign \new_Sorter100|3379_  = \new_Sorter100|3279_  & \new_Sorter100|3280_ ;
  assign \new_Sorter100|3380_  = \new_Sorter100|3279_  | \new_Sorter100|3280_ ;
  assign \new_Sorter100|3381_  = \new_Sorter100|3281_  & \new_Sorter100|3282_ ;
  assign \new_Sorter100|3382_  = \new_Sorter100|3281_  | \new_Sorter100|3282_ ;
  assign \new_Sorter100|3383_  = \new_Sorter100|3283_  & \new_Sorter100|3284_ ;
  assign \new_Sorter100|3384_  = \new_Sorter100|3283_  | \new_Sorter100|3284_ ;
  assign \new_Sorter100|3385_  = \new_Sorter100|3285_  & \new_Sorter100|3286_ ;
  assign \new_Sorter100|3386_  = \new_Sorter100|3285_  | \new_Sorter100|3286_ ;
  assign \new_Sorter100|3387_  = \new_Sorter100|3287_  & \new_Sorter100|3288_ ;
  assign \new_Sorter100|3388_  = \new_Sorter100|3287_  | \new_Sorter100|3288_ ;
  assign \new_Sorter100|3389_  = \new_Sorter100|3289_  & \new_Sorter100|3290_ ;
  assign \new_Sorter100|3390_  = \new_Sorter100|3289_  | \new_Sorter100|3290_ ;
  assign \new_Sorter100|3391_  = \new_Sorter100|3291_  & \new_Sorter100|3292_ ;
  assign \new_Sorter100|3392_  = \new_Sorter100|3291_  | \new_Sorter100|3292_ ;
  assign \new_Sorter100|3393_  = \new_Sorter100|3293_  & \new_Sorter100|3294_ ;
  assign \new_Sorter100|3394_  = \new_Sorter100|3293_  | \new_Sorter100|3294_ ;
  assign \new_Sorter100|3395_  = \new_Sorter100|3295_  & \new_Sorter100|3296_ ;
  assign \new_Sorter100|3396_  = \new_Sorter100|3295_  | \new_Sorter100|3296_ ;
  assign \new_Sorter100|3397_  = \new_Sorter100|3297_  & \new_Sorter100|3298_ ;
  assign \new_Sorter100|3398_  = \new_Sorter100|3297_  | \new_Sorter100|3298_ ;
  assign \new_Sorter100|3400_  = \new_Sorter100|3300_  & \new_Sorter100|3301_ ;
  assign \new_Sorter100|3401_  = \new_Sorter100|3300_  | \new_Sorter100|3301_ ;
  assign \new_Sorter100|3402_  = \new_Sorter100|3302_  & \new_Sorter100|3303_ ;
  assign \new_Sorter100|3403_  = \new_Sorter100|3302_  | \new_Sorter100|3303_ ;
  assign \new_Sorter100|3404_  = \new_Sorter100|3304_  & \new_Sorter100|3305_ ;
  assign \new_Sorter100|3405_  = \new_Sorter100|3304_  | \new_Sorter100|3305_ ;
  assign \new_Sorter100|3406_  = \new_Sorter100|3306_  & \new_Sorter100|3307_ ;
  assign \new_Sorter100|3407_  = \new_Sorter100|3306_  | \new_Sorter100|3307_ ;
  assign \new_Sorter100|3408_  = \new_Sorter100|3308_  & \new_Sorter100|3309_ ;
  assign \new_Sorter100|3409_  = \new_Sorter100|3308_  | \new_Sorter100|3309_ ;
  assign \new_Sorter100|3410_  = \new_Sorter100|3310_  & \new_Sorter100|3311_ ;
  assign \new_Sorter100|3411_  = \new_Sorter100|3310_  | \new_Sorter100|3311_ ;
  assign \new_Sorter100|3412_  = \new_Sorter100|3312_  & \new_Sorter100|3313_ ;
  assign \new_Sorter100|3413_  = \new_Sorter100|3312_  | \new_Sorter100|3313_ ;
  assign \new_Sorter100|3414_  = \new_Sorter100|3314_  & \new_Sorter100|3315_ ;
  assign \new_Sorter100|3415_  = \new_Sorter100|3314_  | \new_Sorter100|3315_ ;
  assign \new_Sorter100|3416_  = \new_Sorter100|3316_  & \new_Sorter100|3317_ ;
  assign \new_Sorter100|3417_  = \new_Sorter100|3316_  | \new_Sorter100|3317_ ;
  assign \new_Sorter100|3418_  = \new_Sorter100|3318_  & \new_Sorter100|3319_ ;
  assign \new_Sorter100|3419_  = \new_Sorter100|3318_  | \new_Sorter100|3319_ ;
  assign \new_Sorter100|3420_  = \new_Sorter100|3320_  & \new_Sorter100|3321_ ;
  assign \new_Sorter100|3421_  = \new_Sorter100|3320_  | \new_Sorter100|3321_ ;
  assign \new_Sorter100|3422_  = \new_Sorter100|3322_  & \new_Sorter100|3323_ ;
  assign \new_Sorter100|3423_  = \new_Sorter100|3322_  | \new_Sorter100|3323_ ;
  assign \new_Sorter100|3424_  = \new_Sorter100|3324_  & \new_Sorter100|3325_ ;
  assign \new_Sorter100|3425_  = \new_Sorter100|3324_  | \new_Sorter100|3325_ ;
  assign \new_Sorter100|3426_  = \new_Sorter100|3326_  & \new_Sorter100|3327_ ;
  assign \new_Sorter100|3427_  = \new_Sorter100|3326_  | \new_Sorter100|3327_ ;
  assign \new_Sorter100|3428_  = \new_Sorter100|3328_  & \new_Sorter100|3329_ ;
  assign \new_Sorter100|3429_  = \new_Sorter100|3328_  | \new_Sorter100|3329_ ;
  assign \new_Sorter100|3430_  = \new_Sorter100|3330_  & \new_Sorter100|3331_ ;
  assign \new_Sorter100|3431_  = \new_Sorter100|3330_  | \new_Sorter100|3331_ ;
  assign \new_Sorter100|3432_  = \new_Sorter100|3332_  & \new_Sorter100|3333_ ;
  assign \new_Sorter100|3433_  = \new_Sorter100|3332_  | \new_Sorter100|3333_ ;
  assign \new_Sorter100|3434_  = \new_Sorter100|3334_  & \new_Sorter100|3335_ ;
  assign \new_Sorter100|3435_  = \new_Sorter100|3334_  | \new_Sorter100|3335_ ;
  assign \new_Sorter100|3436_  = \new_Sorter100|3336_  & \new_Sorter100|3337_ ;
  assign \new_Sorter100|3437_  = \new_Sorter100|3336_  | \new_Sorter100|3337_ ;
  assign \new_Sorter100|3438_  = \new_Sorter100|3338_  & \new_Sorter100|3339_ ;
  assign \new_Sorter100|3439_  = \new_Sorter100|3338_  | \new_Sorter100|3339_ ;
  assign \new_Sorter100|3440_  = \new_Sorter100|3340_  & \new_Sorter100|3341_ ;
  assign \new_Sorter100|3441_  = \new_Sorter100|3340_  | \new_Sorter100|3341_ ;
  assign \new_Sorter100|3442_  = \new_Sorter100|3342_  & \new_Sorter100|3343_ ;
  assign \new_Sorter100|3443_  = \new_Sorter100|3342_  | \new_Sorter100|3343_ ;
  assign \new_Sorter100|3444_  = \new_Sorter100|3344_  & \new_Sorter100|3345_ ;
  assign \new_Sorter100|3445_  = \new_Sorter100|3344_  | \new_Sorter100|3345_ ;
  assign \new_Sorter100|3446_  = \new_Sorter100|3346_  & \new_Sorter100|3347_ ;
  assign \new_Sorter100|3447_  = \new_Sorter100|3346_  | \new_Sorter100|3347_ ;
  assign \new_Sorter100|3448_  = \new_Sorter100|3348_  & \new_Sorter100|3349_ ;
  assign \new_Sorter100|3449_  = \new_Sorter100|3348_  | \new_Sorter100|3349_ ;
  assign \new_Sorter100|3450_  = \new_Sorter100|3350_  & \new_Sorter100|3351_ ;
  assign \new_Sorter100|3451_  = \new_Sorter100|3350_  | \new_Sorter100|3351_ ;
  assign \new_Sorter100|3452_  = \new_Sorter100|3352_  & \new_Sorter100|3353_ ;
  assign \new_Sorter100|3453_  = \new_Sorter100|3352_  | \new_Sorter100|3353_ ;
  assign \new_Sorter100|3454_  = \new_Sorter100|3354_  & \new_Sorter100|3355_ ;
  assign \new_Sorter100|3455_  = \new_Sorter100|3354_  | \new_Sorter100|3355_ ;
  assign \new_Sorter100|3456_  = \new_Sorter100|3356_  & \new_Sorter100|3357_ ;
  assign \new_Sorter100|3457_  = \new_Sorter100|3356_  | \new_Sorter100|3357_ ;
  assign \new_Sorter100|3458_  = \new_Sorter100|3358_  & \new_Sorter100|3359_ ;
  assign \new_Sorter100|3459_  = \new_Sorter100|3358_  | \new_Sorter100|3359_ ;
  assign \new_Sorter100|3460_  = \new_Sorter100|3360_  & \new_Sorter100|3361_ ;
  assign \new_Sorter100|3461_  = \new_Sorter100|3360_  | \new_Sorter100|3361_ ;
  assign \new_Sorter100|3462_  = \new_Sorter100|3362_  & \new_Sorter100|3363_ ;
  assign \new_Sorter100|3463_  = \new_Sorter100|3362_  | \new_Sorter100|3363_ ;
  assign \new_Sorter100|3464_  = \new_Sorter100|3364_  & \new_Sorter100|3365_ ;
  assign \new_Sorter100|3465_  = \new_Sorter100|3364_  | \new_Sorter100|3365_ ;
  assign \new_Sorter100|3466_  = \new_Sorter100|3366_  & \new_Sorter100|3367_ ;
  assign \new_Sorter100|3467_  = \new_Sorter100|3366_  | \new_Sorter100|3367_ ;
  assign \new_Sorter100|3468_  = \new_Sorter100|3368_  & \new_Sorter100|3369_ ;
  assign \new_Sorter100|3469_  = \new_Sorter100|3368_  | \new_Sorter100|3369_ ;
  assign \new_Sorter100|3470_  = \new_Sorter100|3370_  & \new_Sorter100|3371_ ;
  assign \new_Sorter100|3471_  = \new_Sorter100|3370_  | \new_Sorter100|3371_ ;
  assign \new_Sorter100|3472_  = \new_Sorter100|3372_  & \new_Sorter100|3373_ ;
  assign \new_Sorter100|3473_  = \new_Sorter100|3372_  | \new_Sorter100|3373_ ;
  assign \new_Sorter100|3474_  = \new_Sorter100|3374_  & \new_Sorter100|3375_ ;
  assign \new_Sorter100|3475_  = \new_Sorter100|3374_  | \new_Sorter100|3375_ ;
  assign \new_Sorter100|3476_  = \new_Sorter100|3376_  & \new_Sorter100|3377_ ;
  assign \new_Sorter100|3477_  = \new_Sorter100|3376_  | \new_Sorter100|3377_ ;
  assign \new_Sorter100|3478_  = \new_Sorter100|3378_  & \new_Sorter100|3379_ ;
  assign \new_Sorter100|3479_  = \new_Sorter100|3378_  | \new_Sorter100|3379_ ;
  assign \new_Sorter100|3480_  = \new_Sorter100|3380_  & \new_Sorter100|3381_ ;
  assign \new_Sorter100|3481_  = \new_Sorter100|3380_  | \new_Sorter100|3381_ ;
  assign \new_Sorter100|3482_  = \new_Sorter100|3382_  & \new_Sorter100|3383_ ;
  assign \new_Sorter100|3483_  = \new_Sorter100|3382_  | \new_Sorter100|3383_ ;
  assign \new_Sorter100|3484_  = \new_Sorter100|3384_  & \new_Sorter100|3385_ ;
  assign \new_Sorter100|3485_  = \new_Sorter100|3384_  | \new_Sorter100|3385_ ;
  assign \new_Sorter100|3486_  = \new_Sorter100|3386_  & \new_Sorter100|3387_ ;
  assign \new_Sorter100|3487_  = \new_Sorter100|3386_  | \new_Sorter100|3387_ ;
  assign \new_Sorter100|3488_  = \new_Sorter100|3388_  & \new_Sorter100|3389_ ;
  assign \new_Sorter100|3489_  = \new_Sorter100|3388_  | \new_Sorter100|3389_ ;
  assign \new_Sorter100|3490_  = \new_Sorter100|3390_  & \new_Sorter100|3391_ ;
  assign \new_Sorter100|3491_  = \new_Sorter100|3390_  | \new_Sorter100|3391_ ;
  assign \new_Sorter100|3492_  = \new_Sorter100|3392_  & \new_Sorter100|3393_ ;
  assign \new_Sorter100|3493_  = \new_Sorter100|3392_  | \new_Sorter100|3393_ ;
  assign \new_Sorter100|3494_  = \new_Sorter100|3394_  & \new_Sorter100|3395_ ;
  assign \new_Sorter100|3495_  = \new_Sorter100|3394_  | \new_Sorter100|3395_ ;
  assign \new_Sorter100|3496_  = \new_Sorter100|3396_  & \new_Sorter100|3397_ ;
  assign \new_Sorter100|3497_  = \new_Sorter100|3396_  | \new_Sorter100|3397_ ;
  assign \new_Sorter100|3498_  = \new_Sorter100|3398_  & \new_Sorter100|3399_ ;
  assign \new_Sorter100|3499_  = \new_Sorter100|3398_  | \new_Sorter100|3399_ ;
  assign \new_Sorter100|3500_  = \new_Sorter100|3400_ ;
  assign \new_Sorter100|3599_  = \new_Sorter100|3499_ ;
  assign \new_Sorter100|3501_  = \new_Sorter100|3401_  & \new_Sorter100|3402_ ;
  assign \new_Sorter100|3502_  = \new_Sorter100|3401_  | \new_Sorter100|3402_ ;
  assign \new_Sorter100|3503_  = \new_Sorter100|3403_  & \new_Sorter100|3404_ ;
  assign \new_Sorter100|3504_  = \new_Sorter100|3403_  | \new_Sorter100|3404_ ;
  assign \new_Sorter100|3505_  = \new_Sorter100|3405_  & \new_Sorter100|3406_ ;
  assign \new_Sorter100|3506_  = \new_Sorter100|3405_  | \new_Sorter100|3406_ ;
  assign \new_Sorter100|3507_  = \new_Sorter100|3407_  & \new_Sorter100|3408_ ;
  assign \new_Sorter100|3508_  = \new_Sorter100|3407_  | \new_Sorter100|3408_ ;
  assign \new_Sorter100|3509_  = \new_Sorter100|3409_  & \new_Sorter100|3410_ ;
  assign \new_Sorter100|3510_  = \new_Sorter100|3409_  | \new_Sorter100|3410_ ;
  assign \new_Sorter100|3511_  = \new_Sorter100|3411_  & \new_Sorter100|3412_ ;
  assign \new_Sorter100|3512_  = \new_Sorter100|3411_  | \new_Sorter100|3412_ ;
  assign \new_Sorter100|3513_  = \new_Sorter100|3413_  & \new_Sorter100|3414_ ;
  assign \new_Sorter100|3514_  = \new_Sorter100|3413_  | \new_Sorter100|3414_ ;
  assign \new_Sorter100|3515_  = \new_Sorter100|3415_  & \new_Sorter100|3416_ ;
  assign \new_Sorter100|3516_  = \new_Sorter100|3415_  | \new_Sorter100|3416_ ;
  assign \new_Sorter100|3517_  = \new_Sorter100|3417_  & \new_Sorter100|3418_ ;
  assign \new_Sorter100|3518_  = \new_Sorter100|3417_  | \new_Sorter100|3418_ ;
  assign \new_Sorter100|3519_  = \new_Sorter100|3419_  & \new_Sorter100|3420_ ;
  assign \new_Sorter100|3520_  = \new_Sorter100|3419_  | \new_Sorter100|3420_ ;
  assign \new_Sorter100|3521_  = \new_Sorter100|3421_  & \new_Sorter100|3422_ ;
  assign \new_Sorter100|3522_  = \new_Sorter100|3421_  | \new_Sorter100|3422_ ;
  assign \new_Sorter100|3523_  = \new_Sorter100|3423_  & \new_Sorter100|3424_ ;
  assign \new_Sorter100|3524_  = \new_Sorter100|3423_  | \new_Sorter100|3424_ ;
  assign \new_Sorter100|3525_  = \new_Sorter100|3425_  & \new_Sorter100|3426_ ;
  assign \new_Sorter100|3526_  = \new_Sorter100|3425_  | \new_Sorter100|3426_ ;
  assign \new_Sorter100|3527_  = \new_Sorter100|3427_  & \new_Sorter100|3428_ ;
  assign \new_Sorter100|3528_  = \new_Sorter100|3427_  | \new_Sorter100|3428_ ;
  assign \new_Sorter100|3529_  = \new_Sorter100|3429_  & \new_Sorter100|3430_ ;
  assign \new_Sorter100|3530_  = \new_Sorter100|3429_  | \new_Sorter100|3430_ ;
  assign \new_Sorter100|3531_  = \new_Sorter100|3431_  & \new_Sorter100|3432_ ;
  assign \new_Sorter100|3532_  = \new_Sorter100|3431_  | \new_Sorter100|3432_ ;
  assign \new_Sorter100|3533_  = \new_Sorter100|3433_  & \new_Sorter100|3434_ ;
  assign \new_Sorter100|3534_  = \new_Sorter100|3433_  | \new_Sorter100|3434_ ;
  assign \new_Sorter100|3535_  = \new_Sorter100|3435_  & \new_Sorter100|3436_ ;
  assign \new_Sorter100|3536_  = \new_Sorter100|3435_  | \new_Sorter100|3436_ ;
  assign \new_Sorter100|3537_  = \new_Sorter100|3437_  & \new_Sorter100|3438_ ;
  assign \new_Sorter100|3538_  = \new_Sorter100|3437_  | \new_Sorter100|3438_ ;
  assign \new_Sorter100|3539_  = \new_Sorter100|3439_  & \new_Sorter100|3440_ ;
  assign \new_Sorter100|3540_  = \new_Sorter100|3439_  | \new_Sorter100|3440_ ;
  assign \new_Sorter100|3541_  = \new_Sorter100|3441_  & \new_Sorter100|3442_ ;
  assign \new_Sorter100|3542_  = \new_Sorter100|3441_  | \new_Sorter100|3442_ ;
  assign \new_Sorter100|3543_  = \new_Sorter100|3443_  & \new_Sorter100|3444_ ;
  assign \new_Sorter100|3544_  = \new_Sorter100|3443_  | \new_Sorter100|3444_ ;
  assign \new_Sorter100|3545_  = \new_Sorter100|3445_  & \new_Sorter100|3446_ ;
  assign \new_Sorter100|3546_  = \new_Sorter100|3445_  | \new_Sorter100|3446_ ;
  assign \new_Sorter100|3547_  = \new_Sorter100|3447_  & \new_Sorter100|3448_ ;
  assign \new_Sorter100|3548_  = \new_Sorter100|3447_  | \new_Sorter100|3448_ ;
  assign \new_Sorter100|3549_  = \new_Sorter100|3449_  & \new_Sorter100|3450_ ;
  assign \new_Sorter100|3550_  = \new_Sorter100|3449_  | \new_Sorter100|3450_ ;
  assign \new_Sorter100|3551_  = \new_Sorter100|3451_  & \new_Sorter100|3452_ ;
  assign \new_Sorter100|3552_  = \new_Sorter100|3451_  | \new_Sorter100|3452_ ;
  assign \new_Sorter100|3553_  = \new_Sorter100|3453_  & \new_Sorter100|3454_ ;
  assign \new_Sorter100|3554_  = \new_Sorter100|3453_  | \new_Sorter100|3454_ ;
  assign \new_Sorter100|3555_  = \new_Sorter100|3455_  & \new_Sorter100|3456_ ;
  assign \new_Sorter100|3556_  = \new_Sorter100|3455_  | \new_Sorter100|3456_ ;
  assign \new_Sorter100|3557_  = \new_Sorter100|3457_  & \new_Sorter100|3458_ ;
  assign \new_Sorter100|3558_  = \new_Sorter100|3457_  | \new_Sorter100|3458_ ;
  assign \new_Sorter100|3559_  = \new_Sorter100|3459_  & \new_Sorter100|3460_ ;
  assign \new_Sorter100|3560_  = \new_Sorter100|3459_  | \new_Sorter100|3460_ ;
  assign \new_Sorter100|3561_  = \new_Sorter100|3461_  & \new_Sorter100|3462_ ;
  assign \new_Sorter100|3562_  = \new_Sorter100|3461_  | \new_Sorter100|3462_ ;
  assign \new_Sorter100|3563_  = \new_Sorter100|3463_  & \new_Sorter100|3464_ ;
  assign \new_Sorter100|3564_  = \new_Sorter100|3463_  | \new_Sorter100|3464_ ;
  assign \new_Sorter100|3565_  = \new_Sorter100|3465_  & \new_Sorter100|3466_ ;
  assign \new_Sorter100|3566_  = \new_Sorter100|3465_  | \new_Sorter100|3466_ ;
  assign \new_Sorter100|3567_  = \new_Sorter100|3467_  & \new_Sorter100|3468_ ;
  assign \new_Sorter100|3568_  = \new_Sorter100|3467_  | \new_Sorter100|3468_ ;
  assign \new_Sorter100|3569_  = \new_Sorter100|3469_  & \new_Sorter100|3470_ ;
  assign \new_Sorter100|3570_  = \new_Sorter100|3469_  | \new_Sorter100|3470_ ;
  assign \new_Sorter100|3571_  = \new_Sorter100|3471_  & \new_Sorter100|3472_ ;
  assign \new_Sorter100|3572_  = \new_Sorter100|3471_  | \new_Sorter100|3472_ ;
  assign \new_Sorter100|3573_  = \new_Sorter100|3473_  & \new_Sorter100|3474_ ;
  assign \new_Sorter100|3574_  = \new_Sorter100|3473_  | \new_Sorter100|3474_ ;
  assign \new_Sorter100|3575_  = \new_Sorter100|3475_  & \new_Sorter100|3476_ ;
  assign \new_Sorter100|3576_  = \new_Sorter100|3475_  | \new_Sorter100|3476_ ;
  assign \new_Sorter100|3577_  = \new_Sorter100|3477_  & \new_Sorter100|3478_ ;
  assign \new_Sorter100|3578_  = \new_Sorter100|3477_  | \new_Sorter100|3478_ ;
  assign \new_Sorter100|3579_  = \new_Sorter100|3479_  & \new_Sorter100|3480_ ;
  assign \new_Sorter100|3580_  = \new_Sorter100|3479_  | \new_Sorter100|3480_ ;
  assign \new_Sorter100|3581_  = \new_Sorter100|3481_  & \new_Sorter100|3482_ ;
  assign \new_Sorter100|3582_  = \new_Sorter100|3481_  | \new_Sorter100|3482_ ;
  assign \new_Sorter100|3583_  = \new_Sorter100|3483_  & \new_Sorter100|3484_ ;
  assign \new_Sorter100|3584_  = \new_Sorter100|3483_  | \new_Sorter100|3484_ ;
  assign \new_Sorter100|3585_  = \new_Sorter100|3485_  & \new_Sorter100|3486_ ;
  assign \new_Sorter100|3586_  = \new_Sorter100|3485_  | \new_Sorter100|3486_ ;
  assign \new_Sorter100|3587_  = \new_Sorter100|3487_  & \new_Sorter100|3488_ ;
  assign \new_Sorter100|3588_  = \new_Sorter100|3487_  | \new_Sorter100|3488_ ;
  assign \new_Sorter100|3589_  = \new_Sorter100|3489_  & \new_Sorter100|3490_ ;
  assign \new_Sorter100|3590_  = \new_Sorter100|3489_  | \new_Sorter100|3490_ ;
  assign \new_Sorter100|3591_  = \new_Sorter100|3491_  & \new_Sorter100|3492_ ;
  assign \new_Sorter100|3592_  = \new_Sorter100|3491_  | \new_Sorter100|3492_ ;
  assign \new_Sorter100|3593_  = \new_Sorter100|3493_  & \new_Sorter100|3494_ ;
  assign \new_Sorter100|3594_  = \new_Sorter100|3493_  | \new_Sorter100|3494_ ;
  assign \new_Sorter100|3595_  = \new_Sorter100|3495_  & \new_Sorter100|3496_ ;
  assign \new_Sorter100|3596_  = \new_Sorter100|3495_  | \new_Sorter100|3496_ ;
  assign \new_Sorter100|3597_  = \new_Sorter100|3497_  & \new_Sorter100|3498_ ;
  assign \new_Sorter100|3598_  = \new_Sorter100|3497_  | \new_Sorter100|3498_ ;
  assign \new_Sorter100|3600_  = \new_Sorter100|3500_  & \new_Sorter100|3501_ ;
  assign \new_Sorter100|3601_  = \new_Sorter100|3500_  | \new_Sorter100|3501_ ;
  assign \new_Sorter100|3602_  = \new_Sorter100|3502_  & \new_Sorter100|3503_ ;
  assign \new_Sorter100|3603_  = \new_Sorter100|3502_  | \new_Sorter100|3503_ ;
  assign \new_Sorter100|3604_  = \new_Sorter100|3504_  & \new_Sorter100|3505_ ;
  assign \new_Sorter100|3605_  = \new_Sorter100|3504_  | \new_Sorter100|3505_ ;
  assign \new_Sorter100|3606_  = \new_Sorter100|3506_  & \new_Sorter100|3507_ ;
  assign \new_Sorter100|3607_  = \new_Sorter100|3506_  | \new_Sorter100|3507_ ;
  assign \new_Sorter100|3608_  = \new_Sorter100|3508_  & \new_Sorter100|3509_ ;
  assign \new_Sorter100|3609_  = \new_Sorter100|3508_  | \new_Sorter100|3509_ ;
  assign \new_Sorter100|3610_  = \new_Sorter100|3510_  & \new_Sorter100|3511_ ;
  assign \new_Sorter100|3611_  = \new_Sorter100|3510_  | \new_Sorter100|3511_ ;
  assign \new_Sorter100|3612_  = \new_Sorter100|3512_  & \new_Sorter100|3513_ ;
  assign \new_Sorter100|3613_  = \new_Sorter100|3512_  | \new_Sorter100|3513_ ;
  assign \new_Sorter100|3614_  = \new_Sorter100|3514_  & \new_Sorter100|3515_ ;
  assign \new_Sorter100|3615_  = \new_Sorter100|3514_  | \new_Sorter100|3515_ ;
  assign \new_Sorter100|3616_  = \new_Sorter100|3516_  & \new_Sorter100|3517_ ;
  assign \new_Sorter100|3617_  = \new_Sorter100|3516_  | \new_Sorter100|3517_ ;
  assign \new_Sorter100|3618_  = \new_Sorter100|3518_  & \new_Sorter100|3519_ ;
  assign \new_Sorter100|3619_  = \new_Sorter100|3518_  | \new_Sorter100|3519_ ;
  assign \new_Sorter100|3620_  = \new_Sorter100|3520_  & \new_Sorter100|3521_ ;
  assign \new_Sorter100|3621_  = \new_Sorter100|3520_  | \new_Sorter100|3521_ ;
  assign \new_Sorter100|3622_  = \new_Sorter100|3522_  & \new_Sorter100|3523_ ;
  assign \new_Sorter100|3623_  = \new_Sorter100|3522_  | \new_Sorter100|3523_ ;
  assign \new_Sorter100|3624_  = \new_Sorter100|3524_  & \new_Sorter100|3525_ ;
  assign \new_Sorter100|3625_  = \new_Sorter100|3524_  | \new_Sorter100|3525_ ;
  assign \new_Sorter100|3626_  = \new_Sorter100|3526_  & \new_Sorter100|3527_ ;
  assign \new_Sorter100|3627_  = \new_Sorter100|3526_  | \new_Sorter100|3527_ ;
  assign \new_Sorter100|3628_  = \new_Sorter100|3528_  & \new_Sorter100|3529_ ;
  assign \new_Sorter100|3629_  = \new_Sorter100|3528_  | \new_Sorter100|3529_ ;
  assign \new_Sorter100|3630_  = \new_Sorter100|3530_  & \new_Sorter100|3531_ ;
  assign \new_Sorter100|3631_  = \new_Sorter100|3530_  | \new_Sorter100|3531_ ;
  assign \new_Sorter100|3632_  = \new_Sorter100|3532_  & \new_Sorter100|3533_ ;
  assign \new_Sorter100|3633_  = \new_Sorter100|3532_  | \new_Sorter100|3533_ ;
  assign \new_Sorter100|3634_  = \new_Sorter100|3534_  & \new_Sorter100|3535_ ;
  assign \new_Sorter100|3635_  = \new_Sorter100|3534_  | \new_Sorter100|3535_ ;
  assign \new_Sorter100|3636_  = \new_Sorter100|3536_  & \new_Sorter100|3537_ ;
  assign \new_Sorter100|3637_  = \new_Sorter100|3536_  | \new_Sorter100|3537_ ;
  assign \new_Sorter100|3638_  = \new_Sorter100|3538_  & \new_Sorter100|3539_ ;
  assign \new_Sorter100|3639_  = \new_Sorter100|3538_  | \new_Sorter100|3539_ ;
  assign \new_Sorter100|3640_  = \new_Sorter100|3540_  & \new_Sorter100|3541_ ;
  assign \new_Sorter100|3641_  = \new_Sorter100|3540_  | \new_Sorter100|3541_ ;
  assign \new_Sorter100|3642_  = \new_Sorter100|3542_  & \new_Sorter100|3543_ ;
  assign \new_Sorter100|3643_  = \new_Sorter100|3542_  | \new_Sorter100|3543_ ;
  assign \new_Sorter100|3644_  = \new_Sorter100|3544_  & \new_Sorter100|3545_ ;
  assign \new_Sorter100|3645_  = \new_Sorter100|3544_  | \new_Sorter100|3545_ ;
  assign \new_Sorter100|3646_  = \new_Sorter100|3546_  & \new_Sorter100|3547_ ;
  assign \new_Sorter100|3647_  = \new_Sorter100|3546_  | \new_Sorter100|3547_ ;
  assign \new_Sorter100|3648_  = \new_Sorter100|3548_  & \new_Sorter100|3549_ ;
  assign \new_Sorter100|3649_  = \new_Sorter100|3548_  | \new_Sorter100|3549_ ;
  assign \new_Sorter100|3650_  = \new_Sorter100|3550_  & \new_Sorter100|3551_ ;
  assign \new_Sorter100|3651_  = \new_Sorter100|3550_  | \new_Sorter100|3551_ ;
  assign \new_Sorter100|3652_  = \new_Sorter100|3552_  & \new_Sorter100|3553_ ;
  assign \new_Sorter100|3653_  = \new_Sorter100|3552_  | \new_Sorter100|3553_ ;
  assign \new_Sorter100|3654_  = \new_Sorter100|3554_  & \new_Sorter100|3555_ ;
  assign \new_Sorter100|3655_  = \new_Sorter100|3554_  | \new_Sorter100|3555_ ;
  assign \new_Sorter100|3656_  = \new_Sorter100|3556_  & \new_Sorter100|3557_ ;
  assign \new_Sorter100|3657_  = \new_Sorter100|3556_  | \new_Sorter100|3557_ ;
  assign \new_Sorter100|3658_  = \new_Sorter100|3558_  & \new_Sorter100|3559_ ;
  assign \new_Sorter100|3659_  = \new_Sorter100|3558_  | \new_Sorter100|3559_ ;
  assign \new_Sorter100|3660_  = \new_Sorter100|3560_  & \new_Sorter100|3561_ ;
  assign \new_Sorter100|3661_  = \new_Sorter100|3560_  | \new_Sorter100|3561_ ;
  assign \new_Sorter100|3662_  = \new_Sorter100|3562_  & \new_Sorter100|3563_ ;
  assign \new_Sorter100|3663_  = \new_Sorter100|3562_  | \new_Sorter100|3563_ ;
  assign \new_Sorter100|3664_  = \new_Sorter100|3564_  & \new_Sorter100|3565_ ;
  assign \new_Sorter100|3665_  = \new_Sorter100|3564_  | \new_Sorter100|3565_ ;
  assign \new_Sorter100|3666_  = \new_Sorter100|3566_  & \new_Sorter100|3567_ ;
  assign \new_Sorter100|3667_  = \new_Sorter100|3566_  | \new_Sorter100|3567_ ;
  assign \new_Sorter100|3668_  = \new_Sorter100|3568_  & \new_Sorter100|3569_ ;
  assign \new_Sorter100|3669_  = \new_Sorter100|3568_  | \new_Sorter100|3569_ ;
  assign \new_Sorter100|3670_  = \new_Sorter100|3570_  & \new_Sorter100|3571_ ;
  assign \new_Sorter100|3671_  = \new_Sorter100|3570_  | \new_Sorter100|3571_ ;
  assign \new_Sorter100|3672_  = \new_Sorter100|3572_  & \new_Sorter100|3573_ ;
  assign \new_Sorter100|3673_  = \new_Sorter100|3572_  | \new_Sorter100|3573_ ;
  assign \new_Sorter100|3674_  = \new_Sorter100|3574_  & \new_Sorter100|3575_ ;
  assign \new_Sorter100|3675_  = \new_Sorter100|3574_  | \new_Sorter100|3575_ ;
  assign \new_Sorter100|3676_  = \new_Sorter100|3576_  & \new_Sorter100|3577_ ;
  assign \new_Sorter100|3677_  = \new_Sorter100|3576_  | \new_Sorter100|3577_ ;
  assign \new_Sorter100|3678_  = \new_Sorter100|3578_  & \new_Sorter100|3579_ ;
  assign \new_Sorter100|3679_  = \new_Sorter100|3578_  | \new_Sorter100|3579_ ;
  assign \new_Sorter100|3680_  = \new_Sorter100|3580_  & \new_Sorter100|3581_ ;
  assign \new_Sorter100|3681_  = \new_Sorter100|3580_  | \new_Sorter100|3581_ ;
  assign \new_Sorter100|3682_  = \new_Sorter100|3582_  & \new_Sorter100|3583_ ;
  assign \new_Sorter100|3683_  = \new_Sorter100|3582_  | \new_Sorter100|3583_ ;
  assign \new_Sorter100|3684_  = \new_Sorter100|3584_  & \new_Sorter100|3585_ ;
  assign \new_Sorter100|3685_  = \new_Sorter100|3584_  | \new_Sorter100|3585_ ;
  assign \new_Sorter100|3686_  = \new_Sorter100|3586_  & \new_Sorter100|3587_ ;
  assign \new_Sorter100|3687_  = \new_Sorter100|3586_  | \new_Sorter100|3587_ ;
  assign \new_Sorter100|3688_  = \new_Sorter100|3588_  & \new_Sorter100|3589_ ;
  assign \new_Sorter100|3689_  = \new_Sorter100|3588_  | \new_Sorter100|3589_ ;
  assign \new_Sorter100|3690_  = \new_Sorter100|3590_  & \new_Sorter100|3591_ ;
  assign \new_Sorter100|3691_  = \new_Sorter100|3590_  | \new_Sorter100|3591_ ;
  assign \new_Sorter100|3692_  = \new_Sorter100|3592_  & \new_Sorter100|3593_ ;
  assign \new_Sorter100|3693_  = \new_Sorter100|3592_  | \new_Sorter100|3593_ ;
  assign \new_Sorter100|3694_  = \new_Sorter100|3594_  & \new_Sorter100|3595_ ;
  assign \new_Sorter100|3695_  = \new_Sorter100|3594_  | \new_Sorter100|3595_ ;
  assign \new_Sorter100|3696_  = \new_Sorter100|3596_  & \new_Sorter100|3597_ ;
  assign \new_Sorter100|3697_  = \new_Sorter100|3596_  | \new_Sorter100|3597_ ;
  assign \new_Sorter100|3698_  = \new_Sorter100|3598_  & \new_Sorter100|3599_ ;
  assign \new_Sorter100|3699_  = \new_Sorter100|3598_  | \new_Sorter100|3599_ ;
  assign \new_Sorter100|3700_  = \new_Sorter100|3600_ ;
  assign \new_Sorter100|3799_  = \new_Sorter100|3699_ ;
  assign \new_Sorter100|3701_  = \new_Sorter100|3601_  & \new_Sorter100|3602_ ;
  assign \new_Sorter100|3702_  = \new_Sorter100|3601_  | \new_Sorter100|3602_ ;
  assign \new_Sorter100|3703_  = \new_Sorter100|3603_  & \new_Sorter100|3604_ ;
  assign \new_Sorter100|3704_  = \new_Sorter100|3603_  | \new_Sorter100|3604_ ;
  assign \new_Sorter100|3705_  = \new_Sorter100|3605_  & \new_Sorter100|3606_ ;
  assign \new_Sorter100|3706_  = \new_Sorter100|3605_  | \new_Sorter100|3606_ ;
  assign \new_Sorter100|3707_  = \new_Sorter100|3607_  & \new_Sorter100|3608_ ;
  assign \new_Sorter100|3708_  = \new_Sorter100|3607_  | \new_Sorter100|3608_ ;
  assign \new_Sorter100|3709_  = \new_Sorter100|3609_  & \new_Sorter100|3610_ ;
  assign \new_Sorter100|3710_  = \new_Sorter100|3609_  | \new_Sorter100|3610_ ;
  assign \new_Sorter100|3711_  = \new_Sorter100|3611_  & \new_Sorter100|3612_ ;
  assign \new_Sorter100|3712_  = \new_Sorter100|3611_  | \new_Sorter100|3612_ ;
  assign \new_Sorter100|3713_  = \new_Sorter100|3613_  & \new_Sorter100|3614_ ;
  assign \new_Sorter100|3714_  = \new_Sorter100|3613_  | \new_Sorter100|3614_ ;
  assign \new_Sorter100|3715_  = \new_Sorter100|3615_  & \new_Sorter100|3616_ ;
  assign \new_Sorter100|3716_  = \new_Sorter100|3615_  | \new_Sorter100|3616_ ;
  assign \new_Sorter100|3717_  = \new_Sorter100|3617_  & \new_Sorter100|3618_ ;
  assign \new_Sorter100|3718_  = \new_Sorter100|3617_  | \new_Sorter100|3618_ ;
  assign \new_Sorter100|3719_  = \new_Sorter100|3619_  & \new_Sorter100|3620_ ;
  assign \new_Sorter100|3720_  = \new_Sorter100|3619_  | \new_Sorter100|3620_ ;
  assign \new_Sorter100|3721_  = \new_Sorter100|3621_  & \new_Sorter100|3622_ ;
  assign \new_Sorter100|3722_  = \new_Sorter100|3621_  | \new_Sorter100|3622_ ;
  assign \new_Sorter100|3723_  = \new_Sorter100|3623_  & \new_Sorter100|3624_ ;
  assign \new_Sorter100|3724_  = \new_Sorter100|3623_  | \new_Sorter100|3624_ ;
  assign \new_Sorter100|3725_  = \new_Sorter100|3625_  & \new_Sorter100|3626_ ;
  assign \new_Sorter100|3726_  = \new_Sorter100|3625_  | \new_Sorter100|3626_ ;
  assign \new_Sorter100|3727_  = \new_Sorter100|3627_  & \new_Sorter100|3628_ ;
  assign \new_Sorter100|3728_  = \new_Sorter100|3627_  | \new_Sorter100|3628_ ;
  assign \new_Sorter100|3729_  = \new_Sorter100|3629_  & \new_Sorter100|3630_ ;
  assign \new_Sorter100|3730_  = \new_Sorter100|3629_  | \new_Sorter100|3630_ ;
  assign \new_Sorter100|3731_  = \new_Sorter100|3631_  & \new_Sorter100|3632_ ;
  assign \new_Sorter100|3732_  = \new_Sorter100|3631_  | \new_Sorter100|3632_ ;
  assign \new_Sorter100|3733_  = \new_Sorter100|3633_  & \new_Sorter100|3634_ ;
  assign \new_Sorter100|3734_  = \new_Sorter100|3633_  | \new_Sorter100|3634_ ;
  assign \new_Sorter100|3735_  = \new_Sorter100|3635_  & \new_Sorter100|3636_ ;
  assign \new_Sorter100|3736_  = \new_Sorter100|3635_  | \new_Sorter100|3636_ ;
  assign \new_Sorter100|3737_  = \new_Sorter100|3637_  & \new_Sorter100|3638_ ;
  assign \new_Sorter100|3738_  = \new_Sorter100|3637_  | \new_Sorter100|3638_ ;
  assign \new_Sorter100|3739_  = \new_Sorter100|3639_  & \new_Sorter100|3640_ ;
  assign \new_Sorter100|3740_  = \new_Sorter100|3639_  | \new_Sorter100|3640_ ;
  assign \new_Sorter100|3741_  = \new_Sorter100|3641_  & \new_Sorter100|3642_ ;
  assign \new_Sorter100|3742_  = \new_Sorter100|3641_  | \new_Sorter100|3642_ ;
  assign \new_Sorter100|3743_  = \new_Sorter100|3643_  & \new_Sorter100|3644_ ;
  assign \new_Sorter100|3744_  = \new_Sorter100|3643_  | \new_Sorter100|3644_ ;
  assign \new_Sorter100|3745_  = \new_Sorter100|3645_  & \new_Sorter100|3646_ ;
  assign \new_Sorter100|3746_  = \new_Sorter100|3645_  | \new_Sorter100|3646_ ;
  assign \new_Sorter100|3747_  = \new_Sorter100|3647_  & \new_Sorter100|3648_ ;
  assign \new_Sorter100|3748_  = \new_Sorter100|3647_  | \new_Sorter100|3648_ ;
  assign \new_Sorter100|3749_  = \new_Sorter100|3649_  & \new_Sorter100|3650_ ;
  assign \new_Sorter100|3750_  = \new_Sorter100|3649_  | \new_Sorter100|3650_ ;
  assign \new_Sorter100|3751_  = \new_Sorter100|3651_  & \new_Sorter100|3652_ ;
  assign \new_Sorter100|3752_  = \new_Sorter100|3651_  | \new_Sorter100|3652_ ;
  assign \new_Sorter100|3753_  = \new_Sorter100|3653_  & \new_Sorter100|3654_ ;
  assign \new_Sorter100|3754_  = \new_Sorter100|3653_  | \new_Sorter100|3654_ ;
  assign \new_Sorter100|3755_  = \new_Sorter100|3655_  & \new_Sorter100|3656_ ;
  assign \new_Sorter100|3756_  = \new_Sorter100|3655_  | \new_Sorter100|3656_ ;
  assign \new_Sorter100|3757_  = \new_Sorter100|3657_  & \new_Sorter100|3658_ ;
  assign \new_Sorter100|3758_  = \new_Sorter100|3657_  | \new_Sorter100|3658_ ;
  assign \new_Sorter100|3759_  = \new_Sorter100|3659_  & \new_Sorter100|3660_ ;
  assign \new_Sorter100|3760_  = \new_Sorter100|3659_  | \new_Sorter100|3660_ ;
  assign \new_Sorter100|3761_  = \new_Sorter100|3661_  & \new_Sorter100|3662_ ;
  assign \new_Sorter100|3762_  = \new_Sorter100|3661_  | \new_Sorter100|3662_ ;
  assign \new_Sorter100|3763_  = \new_Sorter100|3663_  & \new_Sorter100|3664_ ;
  assign \new_Sorter100|3764_  = \new_Sorter100|3663_  | \new_Sorter100|3664_ ;
  assign \new_Sorter100|3765_  = \new_Sorter100|3665_  & \new_Sorter100|3666_ ;
  assign \new_Sorter100|3766_  = \new_Sorter100|3665_  | \new_Sorter100|3666_ ;
  assign \new_Sorter100|3767_  = \new_Sorter100|3667_  & \new_Sorter100|3668_ ;
  assign \new_Sorter100|3768_  = \new_Sorter100|3667_  | \new_Sorter100|3668_ ;
  assign \new_Sorter100|3769_  = \new_Sorter100|3669_  & \new_Sorter100|3670_ ;
  assign \new_Sorter100|3770_  = \new_Sorter100|3669_  | \new_Sorter100|3670_ ;
  assign \new_Sorter100|3771_  = \new_Sorter100|3671_  & \new_Sorter100|3672_ ;
  assign \new_Sorter100|3772_  = \new_Sorter100|3671_  | \new_Sorter100|3672_ ;
  assign \new_Sorter100|3773_  = \new_Sorter100|3673_  & \new_Sorter100|3674_ ;
  assign \new_Sorter100|3774_  = \new_Sorter100|3673_  | \new_Sorter100|3674_ ;
  assign \new_Sorter100|3775_  = \new_Sorter100|3675_  & \new_Sorter100|3676_ ;
  assign \new_Sorter100|3776_  = \new_Sorter100|3675_  | \new_Sorter100|3676_ ;
  assign \new_Sorter100|3777_  = \new_Sorter100|3677_  & \new_Sorter100|3678_ ;
  assign \new_Sorter100|3778_  = \new_Sorter100|3677_  | \new_Sorter100|3678_ ;
  assign \new_Sorter100|3779_  = \new_Sorter100|3679_  & \new_Sorter100|3680_ ;
  assign \new_Sorter100|3780_  = \new_Sorter100|3679_  | \new_Sorter100|3680_ ;
  assign \new_Sorter100|3781_  = \new_Sorter100|3681_  & \new_Sorter100|3682_ ;
  assign \new_Sorter100|3782_  = \new_Sorter100|3681_  | \new_Sorter100|3682_ ;
  assign \new_Sorter100|3783_  = \new_Sorter100|3683_  & \new_Sorter100|3684_ ;
  assign \new_Sorter100|3784_  = \new_Sorter100|3683_  | \new_Sorter100|3684_ ;
  assign \new_Sorter100|3785_  = \new_Sorter100|3685_  & \new_Sorter100|3686_ ;
  assign \new_Sorter100|3786_  = \new_Sorter100|3685_  | \new_Sorter100|3686_ ;
  assign \new_Sorter100|3787_  = \new_Sorter100|3687_  & \new_Sorter100|3688_ ;
  assign \new_Sorter100|3788_  = \new_Sorter100|3687_  | \new_Sorter100|3688_ ;
  assign \new_Sorter100|3789_  = \new_Sorter100|3689_  & \new_Sorter100|3690_ ;
  assign \new_Sorter100|3790_  = \new_Sorter100|3689_  | \new_Sorter100|3690_ ;
  assign \new_Sorter100|3791_  = \new_Sorter100|3691_  & \new_Sorter100|3692_ ;
  assign \new_Sorter100|3792_  = \new_Sorter100|3691_  | \new_Sorter100|3692_ ;
  assign \new_Sorter100|3793_  = \new_Sorter100|3693_  & \new_Sorter100|3694_ ;
  assign \new_Sorter100|3794_  = \new_Sorter100|3693_  | \new_Sorter100|3694_ ;
  assign \new_Sorter100|3795_  = \new_Sorter100|3695_  & \new_Sorter100|3696_ ;
  assign \new_Sorter100|3796_  = \new_Sorter100|3695_  | \new_Sorter100|3696_ ;
  assign \new_Sorter100|3797_  = \new_Sorter100|3697_  & \new_Sorter100|3698_ ;
  assign \new_Sorter100|3798_  = \new_Sorter100|3697_  | \new_Sorter100|3698_ ;
  assign \new_Sorter100|3800_  = \new_Sorter100|3700_  & \new_Sorter100|3701_ ;
  assign \new_Sorter100|3801_  = \new_Sorter100|3700_  | \new_Sorter100|3701_ ;
  assign \new_Sorter100|3802_  = \new_Sorter100|3702_  & \new_Sorter100|3703_ ;
  assign \new_Sorter100|3803_  = \new_Sorter100|3702_  | \new_Sorter100|3703_ ;
  assign \new_Sorter100|3804_  = \new_Sorter100|3704_  & \new_Sorter100|3705_ ;
  assign \new_Sorter100|3805_  = \new_Sorter100|3704_  | \new_Sorter100|3705_ ;
  assign \new_Sorter100|3806_  = \new_Sorter100|3706_  & \new_Sorter100|3707_ ;
  assign \new_Sorter100|3807_  = \new_Sorter100|3706_  | \new_Sorter100|3707_ ;
  assign \new_Sorter100|3808_  = \new_Sorter100|3708_  & \new_Sorter100|3709_ ;
  assign \new_Sorter100|3809_  = \new_Sorter100|3708_  | \new_Sorter100|3709_ ;
  assign \new_Sorter100|3810_  = \new_Sorter100|3710_  & \new_Sorter100|3711_ ;
  assign \new_Sorter100|3811_  = \new_Sorter100|3710_  | \new_Sorter100|3711_ ;
  assign \new_Sorter100|3812_  = \new_Sorter100|3712_  & \new_Sorter100|3713_ ;
  assign \new_Sorter100|3813_  = \new_Sorter100|3712_  | \new_Sorter100|3713_ ;
  assign \new_Sorter100|3814_  = \new_Sorter100|3714_  & \new_Sorter100|3715_ ;
  assign \new_Sorter100|3815_  = \new_Sorter100|3714_  | \new_Sorter100|3715_ ;
  assign \new_Sorter100|3816_  = \new_Sorter100|3716_  & \new_Sorter100|3717_ ;
  assign \new_Sorter100|3817_  = \new_Sorter100|3716_  | \new_Sorter100|3717_ ;
  assign \new_Sorter100|3818_  = \new_Sorter100|3718_  & \new_Sorter100|3719_ ;
  assign \new_Sorter100|3819_  = \new_Sorter100|3718_  | \new_Sorter100|3719_ ;
  assign \new_Sorter100|3820_  = \new_Sorter100|3720_  & \new_Sorter100|3721_ ;
  assign \new_Sorter100|3821_  = \new_Sorter100|3720_  | \new_Sorter100|3721_ ;
  assign \new_Sorter100|3822_  = \new_Sorter100|3722_  & \new_Sorter100|3723_ ;
  assign \new_Sorter100|3823_  = \new_Sorter100|3722_  | \new_Sorter100|3723_ ;
  assign \new_Sorter100|3824_  = \new_Sorter100|3724_  & \new_Sorter100|3725_ ;
  assign \new_Sorter100|3825_  = \new_Sorter100|3724_  | \new_Sorter100|3725_ ;
  assign \new_Sorter100|3826_  = \new_Sorter100|3726_  & \new_Sorter100|3727_ ;
  assign \new_Sorter100|3827_  = \new_Sorter100|3726_  | \new_Sorter100|3727_ ;
  assign \new_Sorter100|3828_  = \new_Sorter100|3728_  & \new_Sorter100|3729_ ;
  assign \new_Sorter100|3829_  = \new_Sorter100|3728_  | \new_Sorter100|3729_ ;
  assign \new_Sorter100|3830_  = \new_Sorter100|3730_  & \new_Sorter100|3731_ ;
  assign \new_Sorter100|3831_  = \new_Sorter100|3730_  | \new_Sorter100|3731_ ;
  assign \new_Sorter100|3832_  = \new_Sorter100|3732_  & \new_Sorter100|3733_ ;
  assign \new_Sorter100|3833_  = \new_Sorter100|3732_  | \new_Sorter100|3733_ ;
  assign \new_Sorter100|3834_  = \new_Sorter100|3734_  & \new_Sorter100|3735_ ;
  assign \new_Sorter100|3835_  = \new_Sorter100|3734_  | \new_Sorter100|3735_ ;
  assign \new_Sorter100|3836_  = \new_Sorter100|3736_  & \new_Sorter100|3737_ ;
  assign \new_Sorter100|3837_  = \new_Sorter100|3736_  | \new_Sorter100|3737_ ;
  assign \new_Sorter100|3838_  = \new_Sorter100|3738_  & \new_Sorter100|3739_ ;
  assign \new_Sorter100|3839_  = \new_Sorter100|3738_  | \new_Sorter100|3739_ ;
  assign \new_Sorter100|3840_  = \new_Sorter100|3740_  & \new_Sorter100|3741_ ;
  assign \new_Sorter100|3841_  = \new_Sorter100|3740_  | \new_Sorter100|3741_ ;
  assign \new_Sorter100|3842_  = \new_Sorter100|3742_  & \new_Sorter100|3743_ ;
  assign \new_Sorter100|3843_  = \new_Sorter100|3742_  | \new_Sorter100|3743_ ;
  assign \new_Sorter100|3844_  = \new_Sorter100|3744_  & \new_Sorter100|3745_ ;
  assign \new_Sorter100|3845_  = \new_Sorter100|3744_  | \new_Sorter100|3745_ ;
  assign \new_Sorter100|3846_  = \new_Sorter100|3746_  & \new_Sorter100|3747_ ;
  assign \new_Sorter100|3847_  = \new_Sorter100|3746_  | \new_Sorter100|3747_ ;
  assign \new_Sorter100|3848_  = \new_Sorter100|3748_  & \new_Sorter100|3749_ ;
  assign \new_Sorter100|3849_  = \new_Sorter100|3748_  | \new_Sorter100|3749_ ;
  assign \new_Sorter100|3850_  = \new_Sorter100|3750_  & \new_Sorter100|3751_ ;
  assign \new_Sorter100|3851_  = \new_Sorter100|3750_  | \new_Sorter100|3751_ ;
  assign \new_Sorter100|3852_  = \new_Sorter100|3752_  & \new_Sorter100|3753_ ;
  assign \new_Sorter100|3853_  = \new_Sorter100|3752_  | \new_Sorter100|3753_ ;
  assign \new_Sorter100|3854_  = \new_Sorter100|3754_  & \new_Sorter100|3755_ ;
  assign \new_Sorter100|3855_  = \new_Sorter100|3754_  | \new_Sorter100|3755_ ;
  assign \new_Sorter100|3856_  = \new_Sorter100|3756_  & \new_Sorter100|3757_ ;
  assign \new_Sorter100|3857_  = \new_Sorter100|3756_  | \new_Sorter100|3757_ ;
  assign \new_Sorter100|3858_  = \new_Sorter100|3758_  & \new_Sorter100|3759_ ;
  assign \new_Sorter100|3859_  = \new_Sorter100|3758_  | \new_Sorter100|3759_ ;
  assign \new_Sorter100|3860_  = \new_Sorter100|3760_  & \new_Sorter100|3761_ ;
  assign \new_Sorter100|3861_  = \new_Sorter100|3760_  | \new_Sorter100|3761_ ;
  assign \new_Sorter100|3862_  = \new_Sorter100|3762_  & \new_Sorter100|3763_ ;
  assign \new_Sorter100|3863_  = \new_Sorter100|3762_  | \new_Sorter100|3763_ ;
  assign \new_Sorter100|3864_  = \new_Sorter100|3764_  & \new_Sorter100|3765_ ;
  assign \new_Sorter100|3865_  = \new_Sorter100|3764_  | \new_Sorter100|3765_ ;
  assign \new_Sorter100|3866_  = \new_Sorter100|3766_  & \new_Sorter100|3767_ ;
  assign \new_Sorter100|3867_  = \new_Sorter100|3766_  | \new_Sorter100|3767_ ;
  assign \new_Sorter100|3868_  = \new_Sorter100|3768_  & \new_Sorter100|3769_ ;
  assign \new_Sorter100|3869_  = \new_Sorter100|3768_  | \new_Sorter100|3769_ ;
  assign \new_Sorter100|3870_  = \new_Sorter100|3770_  & \new_Sorter100|3771_ ;
  assign \new_Sorter100|3871_  = \new_Sorter100|3770_  | \new_Sorter100|3771_ ;
  assign \new_Sorter100|3872_  = \new_Sorter100|3772_  & \new_Sorter100|3773_ ;
  assign \new_Sorter100|3873_  = \new_Sorter100|3772_  | \new_Sorter100|3773_ ;
  assign \new_Sorter100|3874_  = \new_Sorter100|3774_  & \new_Sorter100|3775_ ;
  assign \new_Sorter100|3875_  = \new_Sorter100|3774_  | \new_Sorter100|3775_ ;
  assign \new_Sorter100|3876_  = \new_Sorter100|3776_  & \new_Sorter100|3777_ ;
  assign \new_Sorter100|3877_  = \new_Sorter100|3776_  | \new_Sorter100|3777_ ;
  assign \new_Sorter100|3878_  = \new_Sorter100|3778_  & \new_Sorter100|3779_ ;
  assign \new_Sorter100|3879_  = \new_Sorter100|3778_  | \new_Sorter100|3779_ ;
  assign \new_Sorter100|3880_  = \new_Sorter100|3780_  & \new_Sorter100|3781_ ;
  assign \new_Sorter100|3881_  = \new_Sorter100|3780_  | \new_Sorter100|3781_ ;
  assign \new_Sorter100|3882_  = \new_Sorter100|3782_  & \new_Sorter100|3783_ ;
  assign \new_Sorter100|3883_  = \new_Sorter100|3782_  | \new_Sorter100|3783_ ;
  assign \new_Sorter100|3884_  = \new_Sorter100|3784_  & \new_Sorter100|3785_ ;
  assign \new_Sorter100|3885_  = \new_Sorter100|3784_  | \new_Sorter100|3785_ ;
  assign \new_Sorter100|3886_  = \new_Sorter100|3786_  & \new_Sorter100|3787_ ;
  assign \new_Sorter100|3887_  = \new_Sorter100|3786_  | \new_Sorter100|3787_ ;
  assign \new_Sorter100|3888_  = \new_Sorter100|3788_  & \new_Sorter100|3789_ ;
  assign \new_Sorter100|3889_  = \new_Sorter100|3788_  | \new_Sorter100|3789_ ;
  assign \new_Sorter100|3890_  = \new_Sorter100|3790_  & \new_Sorter100|3791_ ;
  assign \new_Sorter100|3891_  = \new_Sorter100|3790_  | \new_Sorter100|3791_ ;
  assign \new_Sorter100|3892_  = \new_Sorter100|3792_  & \new_Sorter100|3793_ ;
  assign \new_Sorter100|3893_  = \new_Sorter100|3792_  | \new_Sorter100|3793_ ;
  assign \new_Sorter100|3894_  = \new_Sorter100|3794_  & \new_Sorter100|3795_ ;
  assign \new_Sorter100|3895_  = \new_Sorter100|3794_  | \new_Sorter100|3795_ ;
  assign \new_Sorter100|3896_  = \new_Sorter100|3796_  & \new_Sorter100|3797_ ;
  assign \new_Sorter100|3897_  = \new_Sorter100|3796_  | \new_Sorter100|3797_ ;
  assign \new_Sorter100|3898_  = \new_Sorter100|3798_  & \new_Sorter100|3799_ ;
  assign \new_Sorter100|3899_  = \new_Sorter100|3798_  | \new_Sorter100|3799_ ;
  assign \new_Sorter100|3900_  = \new_Sorter100|3800_ ;
  assign \new_Sorter100|3999_  = \new_Sorter100|3899_ ;
  assign \new_Sorter100|3901_  = \new_Sorter100|3801_  & \new_Sorter100|3802_ ;
  assign \new_Sorter100|3902_  = \new_Sorter100|3801_  | \new_Sorter100|3802_ ;
  assign \new_Sorter100|3903_  = \new_Sorter100|3803_  & \new_Sorter100|3804_ ;
  assign \new_Sorter100|3904_  = \new_Sorter100|3803_  | \new_Sorter100|3804_ ;
  assign \new_Sorter100|3905_  = \new_Sorter100|3805_  & \new_Sorter100|3806_ ;
  assign \new_Sorter100|3906_  = \new_Sorter100|3805_  | \new_Sorter100|3806_ ;
  assign \new_Sorter100|3907_  = \new_Sorter100|3807_  & \new_Sorter100|3808_ ;
  assign \new_Sorter100|3908_  = \new_Sorter100|3807_  | \new_Sorter100|3808_ ;
  assign \new_Sorter100|3909_  = \new_Sorter100|3809_  & \new_Sorter100|3810_ ;
  assign \new_Sorter100|3910_  = \new_Sorter100|3809_  | \new_Sorter100|3810_ ;
  assign \new_Sorter100|3911_  = \new_Sorter100|3811_  & \new_Sorter100|3812_ ;
  assign \new_Sorter100|3912_  = \new_Sorter100|3811_  | \new_Sorter100|3812_ ;
  assign \new_Sorter100|3913_  = \new_Sorter100|3813_  & \new_Sorter100|3814_ ;
  assign \new_Sorter100|3914_  = \new_Sorter100|3813_  | \new_Sorter100|3814_ ;
  assign \new_Sorter100|3915_  = \new_Sorter100|3815_  & \new_Sorter100|3816_ ;
  assign \new_Sorter100|3916_  = \new_Sorter100|3815_  | \new_Sorter100|3816_ ;
  assign \new_Sorter100|3917_  = \new_Sorter100|3817_  & \new_Sorter100|3818_ ;
  assign \new_Sorter100|3918_  = \new_Sorter100|3817_  | \new_Sorter100|3818_ ;
  assign \new_Sorter100|3919_  = \new_Sorter100|3819_  & \new_Sorter100|3820_ ;
  assign \new_Sorter100|3920_  = \new_Sorter100|3819_  | \new_Sorter100|3820_ ;
  assign \new_Sorter100|3921_  = \new_Sorter100|3821_  & \new_Sorter100|3822_ ;
  assign \new_Sorter100|3922_  = \new_Sorter100|3821_  | \new_Sorter100|3822_ ;
  assign \new_Sorter100|3923_  = \new_Sorter100|3823_  & \new_Sorter100|3824_ ;
  assign \new_Sorter100|3924_  = \new_Sorter100|3823_  | \new_Sorter100|3824_ ;
  assign \new_Sorter100|3925_  = \new_Sorter100|3825_  & \new_Sorter100|3826_ ;
  assign \new_Sorter100|3926_  = \new_Sorter100|3825_  | \new_Sorter100|3826_ ;
  assign \new_Sorter100|3927_  = \new_Sorter100|3827_  & \new_Sorter100|3828_ ;
  assign \new_Sorter100|3928_  = \new_Sorter100|3827_  | \new_Sorter100|3828_ ;
  assign \new_Sorter100|3929_  = \new_Sorter100|3829_  & \new_Sorter100|3830_ ;
  assign \new_Sorter100|3930_  = \new_Sorter100|3829_  | \new_Sorter100|3830_ ;
  assign \new_Sorter100|3931_  = \new_Sorter100|3831_  & \new_Sorter100|3832_ ;
  assign \new_Sorter100|3932_  = \new_Sorter100|3831_  | \new_Sorter100|3832_ ;
  assign \new_Sorter100|3933_  = \new_Sorter100|3833_  & \new_Sorter100|3834_ ;
  assign \new_Sorter100|3934_  = \new_Sorter100|3833_  | \new_Sorter100|3834_ ;
  assign \new_Sorter100|3935_  = \new_Sorter100|3835_  & \new_Sorter100|3836_ ;
  assign \new_Sorter100|3936_  = \new_Sorter100|3835_  | \new_Sorter100|3836_ ;
  assign \new_Sorter100|3937_  = \new_Sorter100|3837_  & \new_Sorter100|3838_ ;
  assign \new_Sorter100|3938_  = \new_Sorter100|3837_  | \new_Sorter100|3838_ ;
  assign \new_Sorter100|3939_  = \new_Sorter100|3839_  & \new_Sorter100|3840_ ;
  assign \new_Sorter100|3940_  = \new_Sorter100|3839_  | \new_Sorter100|3840_ ;
  assign \new_Sorter100|3941_  = \new_Sorter100|3841_  & \new_Sorter100|3842_ ;
  assign \new_Sorter100|3942_  = \new_Sorter100|3841_  | \new_Sorter100|3842_ ;
  assign \new_Sorter100|3943_  = \new_Sorter100|3843_  & \new_Sorter100|3844_ ;
  assign \new_Sorter100|3944_  = \new_Sorter100|3843_  | \new_Sorter100|3844_ ;
  assign \new_Sorter100|3945_  = \new_Sorter100|3845_  & \new_Sorter100|3846_ ;
  assign \new_Sorter100|3946_  = \new_Sorter100|3845_  | \new_Sorter100|3846_ ;
  assign \new_Sorter100|3947_  = \new_Sorter100|3847_  & \new_Sorter100|3848_ ;
  assign \new_Sorter100|3948_  = \new_Sorter100|3847_  | \new_Sorter100|3848_ ;
  assign \new_Sorter100|3949_  = \new_Sorter100|3849_  & \new_Sorter100|3850_ ;
  assign \new_Sorter100|3950_  = \new_Sorter100|3849_  | \new_Sorter100|3850_ ;
  assign \new_Sorter100|3951_  = \new_Sorter100|3851_  & \new_Sorter100|3852_ ;
  assign \new_Sorter100|3952_  = \new_Sorter100|3851_  | \new_Sorter100|3852_ ;
  assign \new_Sorter100|3953_  = \new_Sorter100|3853_  & \new_Sorter100|3854_ ;
  assign \new_Sorter100|3954_  = \new_Sorter100|3853_  | \new_Sorter100|3854_ ;
  assign \new_Sorter100|3955_  = \new_Sorter100|3855_  & \new_Sorter100|3856_ ;
  assign \new_Sorter100|3956_  = \new_Sorter100|3855_  | \new_Sorter100|3856_ ;
  assign \new_Sorter100|3957_  = \new_Sorter100|3857_  & \new_Sorter100|3858_ ;
  assign \new_Sorter100|3958_  = \new_Sorter100|3857_  | \new_Sorter100|3858_ ;
  assign \new_Sorter100|3959_  = \new_Sorter100|3859_  & \new_Sorter100|3860_ ;
  assign \new_Sorter100|3960_  = \new_Sorter100|3859_  | \new_Sorter100|3860_ ;
  assign \new_Sorter100|3961_  = \new_Sorter100|3861_  & \new_Sorter100|3862_ ;
  assign \new_Sorter100|3962_  = \new_Sorter100|3861_  | \new_Sorter100|3862_ ;
  assign \new_Sorter100|3963_  = \new_Sorter100|3863_  & \new_Sorter100|3864_ ;
  assign \new_Sorter100|3964_  = \new_Sorter100|3863_  | \new_Sorter100|3864_ ;
  assign \new_Sorter100|3965_  = \new_Sorter100|3865_  & \new_Sorter100|3866_ ;
  assign \new_Sorter100|3966_  = \new_Sorter100|3865_  | \new_Sorter100|3866_ ;
  assign \new_Sorter100|3967_  = \new_Sorter100|3867_  & \new_Sorter100|3868_ ;
  assign \new_Sorter100|3968_  = \new_Sorter100|3867_  | \new_Sorter100|3868_ ;
  assign \new_Sorter100|3969_  = \new_Sorter100|3869_  & \new_Sorter100|3870_ ;
  assign \new_Sorter100|3970_  = \new_Sorter100|3869_  | \new_Sorter100|3870_ ;
  assign \new_Sorter100|3971_  = \new_Sorter100|3871_  & \new_Sorter100|3872_ ;
  assign \new_Sorter100|3972_  = \new_Sorter100|3871_  | \new_Sorter100|3872_ ;
  assign \new_Sorter100|3973_  = \new_Sorter100|3873_  & \new_Sorter100|3874_ ;
  assign \new_Sorter100|3974_  = \new_Sorter100|3873_  | \new_Sorter100|3874_ ;
  assign \new_Sorter100|3975_  = \new_Sorter100|3875_  & \new_Sorter100|3876_ ;
  assign \new_Sorter100|3976_  = \new_Sorter100|3875_  | \new_Sorter100|3876_ ;
  assign \new_Sorter100|3977_  = \new_Sorter100|3877_  & \new_Sorter100|3878_ ;
  assign \new_Sorter100|3978_  = \new_Sorter100|3877_  | \new_Sorter100|3878_ ;
  assign \new_Sorter100|3979_  = \new_Sorter100|3879_  & \new_Sorter100|3880_ ;
  assign \new_Sorter100|3980_  = \new_Sorter100|3879_  | \new_Sorter100|3880_ ;
  assign \new_Sorter100|3981_  = \new_Sorter100|3881_  & \new_Sorter100|3882_ ;
  assign \new_Sorter100|3982_  = \new_Sorter100|3881_  | \new_Sorter100|3882_ ;
  assign \new_Sorter100|3983_  = \new_Sorter100|3883_  & \new_Sorter100|3884_ ;
  assign \new_Sorter100|3984_  = \new_Sorter100|3883_  | \new_Sorter100|3884_ ;
  assign \new_Sorter100|3985_  = \new_Sorter100|3885_  & \new_Sorter100|3886_ ;
  assign \new_Sorter100|3986_  = \new_Sorter100|3885_  | \new_Sorter100|3886_ ;
  assign \new_Sorter100|3987_  = \new_Sorter100|3887_  & \new_Sorter100|3888_ ;
  assign \new_Sorter100|3988_  = \new_Sorter100|3887_  | \new_Sorter100|3888_ ;
  assign \new_Sorter100|3989_  = \new_Sorter100|3889_  & \new_Sorter100|3890_ ;
  assign \new_Sorter100|3990_  = \new_Sorter100|3889_  | \new_Sorter100|3890_ ;
  assign \new_Sorter100|3991_  = \new_Sorter100|3891_  & \new_Sorter100|3892_ ;
  assign \new_Sorter100|3992_  = \new_Sorter100|3891_  | \new_Sorter100|3892_ ;
  assign \new_Sorter100|3993_  = \new_Sorter100|3893_  & \new_Sorter100|3894_ ;
  assign \new_Sorter100|3994_  = \new_Sorter100|3893_  | \new_Sorter100|3894_ ;
  assign \new_Sorter100|3995_  = \new_Sorter100|3895_  & \new_Sorter100|3896_ ;
  assign \new_Sorter100|3996_  = \new_Sorter100|3895_  | \new_Sorter100|3896_ ;
  assign \new_Sorter100|3997_  = \new_Sorter100|3897_  & \new_Sorter100|3898_ ;
  assign \new_Sorter100|3998_  = \new_Sorter100|3897_  | \new_Sorter100|3898_ ;
  assign \new_Sorter100|4000_  = \new_Sorter100|3900_  & \new_Sorter100|3901_ ;
  assign \new_Sorter100|4001_  = \new_Sorter100|3900_  | \new_Sorter100|3901_ ;
  assign \new_Sorter100|4002_  = \new_Sorter100|3902_  & \new_Sorter100|3903_ ;
  assign \new_Sorter100|4003_  = \new_Sorter100|3902_  | \new_Sorter100|3903_ ;
  assign \new_Sorter100|4004_  = \new_Sorter100|3904_  & \new_Sorter100|3905_ ;
  assign \new_Sorter100|4005_  = \new_Sorter100|3904_  | \new_Sorter100|3905_ ;
  assign \new_Sorter100|4006_  = \new_Sorter100|3906_  & \new_Sorter100|3907_ ;
  assign \new_Sorter100|4007_  = \new_Sorter100|3906_  | \new_Sorter100|3907_ ;
  assign \new_Sorter100|4008_  = \new_Sorter100|3908_  & \new_Sorter100|3909_ ;
  assign \new_Sorter100|4009_  = \new_Sorter100|3908_  | \new_Sorter100|3909_ ;
  assign \new_Sorter100|4010_  = \new_Sorter100|3910_  & \new_Sorter100|3911_ ;
  assign \new_Sorter100|4011_  = \new_Sorter100|3910_  | \new_Sorter100|3911_ ;
  assign \new_Sorter100|4012_  = \new_Sorter100|3912_  & \new_Sorter100|3913_ ;
  assign \new_Sorter100|4013_  = \new_Sorter100|3912_  | \new_Sorter100|3913_ ;
  assign \new_Sorter100|4014_  = \new_Sorter100|3914_  & \new_Sorter100|3915_ ;
  assign \new_Sorter100|4015_  = \new_Sorter100|3914_  | \new_Sorter100|3915_ ;
  assign \new_Sorter100|4016_  = \new_Sorter100|3916_  & \new_Sorter100|3917_ ;
  assign \new_Sorter100|4017_  = \new_Sorter100|3916_  | \new_Sorter100|3917_ ;
  assign \new_Sorter100|4018_  = \new_Sorter100|3918_  & \new_Sorter100|3919_ ;
  assign \new_Sorter100|4019_  = \new_Sorter100|3918_  | \new_Sorter100|3919_ ;
  assign \new_Sorter100|4020_  = \new_Sorter100|3920_  & \new_Sorter100|3921_ ;
  assign \new_Sorter100|4021_  = \new_Sorter100|3920_  | \new_Sorter100|3921_ ;
  assign \new_Sorter100|4022_  = \new_Sorter100|3922_  & \new_Sorter100|3923_ ;
  assign \new_Sorter100|4023_  = \new_Sorter100|3922_  | \new_Sorter100|3923_ ;
  assign \new_Sorter100|4024_  = \new_Sorter100|3924_  & \new_Sorter100|3925_ ;
  assign \new_Sorter100|4025_  = \new_Sorter100|3924_  | \new_Sorter100|3925_ ;
  assign \new_Sorter100|4026_  = \new_Sorter100|3926_  & \new_Sorter100|3927_ ;
  assign \new_Sorter100|4027_  = \new_Sorter100|3926_  | \new_Sorter100|3927_ ;
  assign \new_Sorter100|4028_  = \new_Sorter100|3928_  & \new_Sorter100|3929_ ;
  assign \new_Sorter100|4029_  = \new_Sorter100|3928_  | \new_Sorter100|3929_ ;
  assign \new_Sorter100|4030_  = \new_Sorter100|3930_  & \new_Sorter100|3931_ ;
  assign \new_Sorter100|4031_  = \new_Sorter100|3930_  | \new_Sorter100|3931_ ;
  assign \new_Sorter100|4032_  = \new_Sorter100|3932_  & \new_Sorter100|3933_ ;
  assign \new_Sorter100|4033_  = \new_Sorter100|3932_  | \new_Sorter100|3933_ ;
  assign \new_Sorter100|4034_  = \new_Sorter100|3934_  & \new_Sorter100|3935_ ;
  assign \new_Sorter100|4035_  = \new_Sorter100|3934_  | \new_Sorter100|3935_ ;
  assign \new_Sorter100|4036_  = \new_Sorter100|3936_  & \new_Sorter100|3937_ ;
  assign \new_Sorter100|4037_  = \new_Sorter100|3936_  | \new_Sorter100|3937_ ;
  assign \new_Sorter100|4038_  = \new_Sorter100|3938_  & \new_Sorter100|3939_ ;
  assign \new_Sorter100|4039_  = \new_Sorter100|3938_  | \new_Sorter100|3939_ ;
  assign \new_Sorter100|4040_  = \new_Sorter100|3940_  & \new_Sorter100|3941_ ;
  assign \new_Sorter100|4041_  = \new_Sorter100|3940_  | \new_Sorter100|3941_ ;
  assign \new_Sorter100|4042_  = \new_Sorter100|3942_  & \new_Sorter100|3943_ ;
  assign \new_Sorter100|4043_  = \new_Sorter100|3942_  | \new_Sorter100|3943_ ;
  assign \new_Sorter100|4044_  = \new_Sorter100|3944_  & \new_Sorter100|3945_ ;
  assign \new_Sorter100|4045_  = \new_Sorter100|3944_  | \new_Sorter100|3945_ ;
  assign \new_Sorter100|4046_  = \new_Sorter100|3946_  & \new_Sorter100|3947_ ;
  assign \new_Sorter100|4047_  = \new_Sorter100|3946_  | \new_Sorter100|3947_ ;
  assign \new_Sorter100|4048_  = \new_Sorter100|3948_  & \new_Sorter100|3949_ ;
  assign \new_Sorter100|4049_  = \new_Sorter100|3948_  | \new_Sorter100|3949_ ;
  assign \new_Sorter100|4050_  = \new_Sorter100|3950_  & \new_Sorter100|3951_ ;
  assign \new_Sorter100|4051_  = \new_Sorter100|3950_  | \new_Sorter100|3951_ ;
  assign \new_Sorter100|4052_  = \new_Sorter100|3952_  & \new_Sorter100|3953_ ;
  assign \new_Sorter100|4053_  = \new_Sorter100|3952_  | \new_Sorter100|3953_ ;
  assign \new_Sorter100|4054_  = \new_Sorter100|3954_  & \new_Sorter100|3955_ ;
  assign \new_Sorter100|4055_  = \new_Sorter100|3954_  | \new_Sorter100|3955_ ;
  assign \new_Sorter100|4056_  = \new_Sorter100|3956_  & \new_Sorter100|3957_ ;
  assign \new_Sorter100|4057_  = \new_Sorter100|3956_  | \new_Sorter100|3957_ ;
  assign \new_Sorter100|4058_  = \new_Sorter100|3958_  & \new_Sorter100|3959_ ;
  assign \new_Sorter100|4059_  = \new_Sorter100|3958_  | \new_Sorter100|3959_ ;
  assign \new_Sorter100|4060_  = \new_Sorter100|3960_  & \new_Sorter100|3961_ ;
  assign \new_Sorter100|4061_  = \new_Sorter100|3960_  | \new_Sorter100|3961_ ;
  assign \new_Sorter100|4062_  = \new_Sorter100|3962_  & \new_Sorter100|3963_ ;
  assign \new_Sorter100|4063_  = \new_Sorter100|3962_  | \new_Sorter100|3963_ ;
  assign \new_Sorter100|4064_  = \new_Sorter100|3964_  & \new_Sorter100|3965_ ;
  assign \new_Sorter100|4065_  = \new_Sorter100|3964_  | \new_Sorter100|3965_ ;
  assign \new_Sorter100|4066_  = \new_Sorter100|3966_  & \new_Sorter100|3967_ ;
  assign \new_Sorter100|4067_  = \new_Sorter100|3966_  | \new_Sorter100|3967_ ;
  assign \new_Sorter100|4068_  = \new_Sorter100|3968_  & \new_Sorter100|3969_ ;
  assign \new_Sorter100|4069_  = \new_Sorter100|3968_  | \new_Sorter100|3969_ ;
  assign \new_Sorter100|4070_  = \new_Sorter100|3970_  & \new_Sorter100|3971_ ;
  assign \new_Sorter100|4071_  = \new_Sorter100|3970_  | \new_Sorter100|3971_ ;
  assign \new_Sorter100|4072_  = \new_Sorter100|3972_  & \new_Sorter100|3973_ ;
  assign \new_Sorter100|4073_  = \new_Sorter100|3972_  | \new_Sorter100|3973_ ;
  assign \new_Sorter100|4074_  = \new_Sorter100|3974_  & \new_Sorter100|3975_ ;
  assign \new_Sorter100|4075_  = \new_Sorter100|3974_  | \new_Sorter100|3975_ ;
  assign \new_Sorter100|4076_  = \new_Sorter100|3976_  & \new_Sorter100|3977_ ;
  assign \new_Sorter100|4077_  = \new_Sorter100|3976_  | \new_Sorter100|3977_ ;
  assign \new_Sorter100|4078_  = \new_Sorter100|3978_  & \new_Sorter100|3979_ ;
  assign \new_Sorter100|4079_  = \new_Sorter100|3978_  | \new_Sorter100|3979_ ;
  assign \new_Sorter100|4080_  = \new_Sorter100|3980_  & \new_Sorter100|3981_ ;
  assign \new_Sorter100|4081_  = \new_Sorter100|3980_  | \new_Sorter100|3981_ ;
  assign \new_Sorter100|4082_  = \new_Sorter100|3982_  & \new_Sorter100|3983_ ;
  assign \new_Sorter100|4083_  = \new_Sorter100|3982_  | \new_Sorter100|3983_ ;
  assign \new_Sorter100|4084_  = \new_Sorter100|3984_  & \new_Sorter100|3985_ ;
  assign \new_Sorter100|4085_  = \new_Sorter100|3984_  | \new_Sorter100|3985_ ;
  assign \new_Sorter100|4086_  = \new_Sorter100|3986_  & \new_Sorter100|3987_ ;
  assign \new_Sorter100|4087_  = \new_Sorter100|3986_  | \new_Sorter100|3987_ ;
  assign \new_Sorter100|4088_  = \new_Sorter100|3988_  & \new_Sorter100|3989_ ;
  assign \new_Sorter100|4089_  = \new_Sorter100|3988_  | \new_Sorter100|3989_ ;
  assign \new_Sorter100|4090_  = \new_Sorter100|3990_  & \new_Sorter100|3991_ ;
  assign \new_Sorter100|4091_  = \new_Sorter100|3990_  | \new_Sorter100|3991_ ;
  assign \new_Sorter100|4092_  = \new_Sorter100|3992_  & \new_Sorter100|3993_ ;
  assign \new_Sorter100|4093_  = \new_Sorter100|3992_  | \new_Sorter100|3993_ ;
  assign \new_Sorter100|4094_  = \new_Sorter100|3994_  & \new_Sorter100|3995_ ;
  assign \new_Sorter100|4095_  = \new_Sorter100|3994_  | \new_Sorter100|3995_ ;
  assign \new_Sorter100|4096_  = \new_Sorter100|3996_  & \new_Sorter100|3997_ ;
  assign \new_Sorter100|4097_  = \new_Sorter100|3996_  | \new_Sorter100|3997_ ;
  assign \new_Sorter100|4098_  = \new_Sorter100|3998_  & \new_Sorter100|3999_ ;
  assign \new_Sorter100|4099_  = \new_Sorter100|3998_  | \new_Sorter100|3999_ ;
  assign \new_Sorter100|4100_  = \new_Sorter100|4000_ ;
  assign \new_Sorter100|4199_  = \new_Sorter100|4099_ ;
  assign \new_Sorter100|4101_  = \new_Sorter100|4001_  & \new_Sorter100|4002_ ;
  assign \new_Sorter100|4102_  = \new_Sorter100|4001_  | \new_Sorter100|4002_ ;
  assign \new_Sorter100|4103_  = \new_Sorter100|4003_  & \new_Sorter100|4004_ ;
  assign \new_Sorter100|4104_  = \new_Sorter100|4003_  | \new_Sorter100|4004_ ;
  assign \new_Sorter100|4105_  = \new_Sorter100|4005_  & \new_Sorter100|4006_ ;
  assign \new_Sorter100|4106_  = \new_Sorter100|4005_  | \new_Sorter100|4006_ ;
  assign \new_Sorter100|4107_  = \new_Sorter100|4007_  & \new_Sorter100|4008_ ;
  assign \new_Sorter100|4108_  = \new_Sorter100|4007_  | \new_Sorter100|4008_ ;
  assign \new_Sorter100|4109_  = \new_Sorter100|4009_  & \new_Sorter100|4010_ ;
  assign \new_Sorter100|4110_  = \new_Sorter100|4009_  | \new_Sorter100|4010_ ;
  assign \new_Sorter100|4111_  = \new_Sorter100|4011_  & \new_Sorter100|4012_ ;
  assign \new_Sorter100|4112_  = \new_Sorter100|4011_  | \new_Sorter100|4012_ ;
  assign \new_Sorter100|4113_  = \new_Sorter100|4013_  & \new_Sorter100|4014_ ;
  assign \new_Sorter100|4114_  = \new_Sorter100|4013_  | \new_Sorter100|4014_ ;
  assign \new_Sorter100|4115_  = \new_Sorter100|4015_  & \new_Sorter100|4016_ ;
  assign \new_Sorter100|4116_  = \new_Sorter100|4015_  | \new_Sorter100|4016_ ;
  assign \new_Sorter100|4117_  = \new_Sorter100|4017_  & \new_Sorter100|4018_ ;
  assign \new_Sorter100|4118_  = \new_Sorter100|4017_  | \new_Sorter100|4018_ ;
  assign \new_Sorter100|4119_  = \new_Sorter100|4019_  & \new_Sorter100|4020_ ;
  assign \new_Sorter100|4120_  = \new_Sorter100|4019_  | \new_Sorter100|4020_ ;
  assign \new_Sorter100|4121_  = \new_Sorter100|4021_  & \new_Sorter100|4022_ ;
  assign \new_Sorter100|4122_  = \new_Sorter100|4021_  | \new_Sorter100|4022_ ;
  assign \new_Sorter100|4123_  = \new_Sorter100|4023_  & \new_Sorter100|4024_ ;
  assign \new_Sorter100|4124_  = \new_Sorter100|4023_  | \new_Sorter100|4024_ ;
  assign \new_Sorter100|4125_  = \new_Sorter100|4025_  & \new_Sorter100|4026_ ;
  assign \new_Sorter100|4126_  = \new_Sorter100|4025_  | \new_Sorter100|4026_ ;
  assign \new_Sorter100|4127_  = \new_Sorter100|4027_  & \new_Sorter100|4028_ ;
  assign \new_Sorter100|4128_  = \new_Sorter100|4027_  | \new_Sorter100|4028_ ;
  assign \new_Sorter100|4129_  = \new_Sorter100|4029_  & \new_Sorter100|4030_ ;
  assign \new_Sorter100|4130_  = \new_Sorter100|4029_  | \new_Sorter100|4030_ ;
  assign \new_Sorter100|4131_  = \new_Sorter100|4031_  & \new_Sorter100|4032_ ;
  assign \new_Sorter100|4132_  = \new_Sorter100|4031_  | \new_Sorter100|4032_ ;
  assign \new_Sorter100|4133_  = \new_Sorter100|4033_  & \new_Sorter100|4034_ ;
  assign \new_Sorter100|4134_  = \new_Sorter100|4033_  | \new_Sorter100|4034_ ;
  assign \new_Sorter100|4135_  = \new_Sorter100|4035_  & \new_Sorter100|4036_ ;
  assign \new_Sorter100|4136_  = \new_Sorter100|4035_  | \new_Sorter100|4036_ ;
  assign \new_Sorter100|4137_  = \new_Sorter100|4037_  & \new_Sorter100|4038_ ;
  assign \new_Sorter100|4138_  = \new_Sorter100|4037_  | \new_Sorter100|4038_ ;
  assign \new_Sorter100|4139_  = \new_Sorter100|4039_  & \new_Sorter100|4040_ ;
  assign \new_Sorter100|4140_  = \new_Sorter100|4039_  | \new_Sorter100|4040_ ;
  assign \new_Sorter100|4141_  = \new_Sorter100|4041_  & \new_Sorter100|4042_ ;
  assign \new_Sorter100|4142_  = \new_Sorter100|4041_  | \new_Sorter100|4042_ ;
  assign \new_Sorter100|4143_  = \new_Sorter100|4043_  & \new_Sorter100|4044_ ;
  assign \new_Sorter100|4144_  = \new_Sorter100|4043_  | \new_Sorter100|4044_ ;
  assign \new_Sorter100|4145_  = \new_Sorter100|4045_  & \new_Sorter100|4046_ ;
  assign \new_Sorter100|4146_  = \new_Sorter100|4045_  | \new_Sorter100|4046_ ;
  assign \new_Sorter100|4147_  = \new_Sorter100|4047_  & \new_Sorter100|4048_ ;
  assign \new_Sorter100|4148_  = \new_Sorter100|4047_  | \new_Sorter100|4048_ ;
  assign \new_Sorter100|4149_  = \new_Sorter100|4049_  & \new_Sorter100|4050_ ;
  assign \new_Sorter100|4150_  = \new_Sorter100|4049_  | \new_Sorter100|4050_ ;
  assign \new_Sorter100|4151_  = \new_Sorter100|4051_  & \new_Sorter100|4052_ ;
  assign \new_Sorter100|4152_  = \new_Sorter100|4051_  | \new_Sorter100|4052_ ;
  assign \new_Sorter100|4153_  = \new_Sorter100|4053_  & \new_Sorter100|4054_ ;
  assign \new_Sorter100|4154_  = \new_Sorter100|4053_  | \new_Sorter100|4054_ ;
  assign \new_Sorter100|4155_  = \new_Sorter100|4055_  & \new_Sorter100|4056_ ;
  assign \new_Sorter100|4156_  = \new_Sorter100|4055_  | \new_Sorter100|4056_ ;
  assign \new_Sorter100|4157_  = \new_Sorter100|4057_  & \new_Sorter100|4058_ ;
  assign \new_Sorter100|4158_  = \new_Sorter100|4057_  | \new_Sorter100|4058_ ;
  assign \new_Sorter100|4159_  = \new_Sorter100|4059_  & \new_Sorter100|4060_ ;
  assign \new_Sorter100|4160_  = \new_Sorter100|4059_  | \new_Sorter100|4060_ ;
  assign \new_Sorter100|4161_  = \new_Sorter100|4061_  & \new_Sorter100|4062_ ;
  assign \new_Sorter100|4162_  = \new_Sorter100|4061_  | \new_Sorter100|4062_ ;
  assign \new_Sorter100|4163_  = \new_Sorter100|4063_  & \new_Sorter100|4064_ ;
  assign \new_Sorter100|4164_  = \new_Sorter100|4063_  | \new_Sorter100|4064_ ;
  assign \new_Sorter100|4165_  = \new_Sorter100|4065_  & \new_Sorter100|4066_ ;
  assign \new_Sorter100|4166_  = \new_Sorter100|4065_  | \new_Sorter100|4066_ ;
  assign \new_Sorter100|4167_  = \new_Sorter100|4067_  & \new_Sorter100|4068_ ;
  assign \new_Sorter100|4168_  = \new_Sorter100|4067_  | \new_Sorter100|4068_ ;
  assign \new_Sorter100|4169_  = \new_Sorter100|4069_  & \new_Sorter100|4070_ ;
  assign \new_Sorter100|4170_  = \new_Sorter100|4069_  | \new_Sorter100|4070_ ;
  assign \new_Sorter100|4171_  = \new_Sorter100|4071_  & \new_Sorter100|4072_ ;
  assign \new_Sorter100|4172_  = \new_Sorter100|4071_  | \new_Sorter100|4072_ ;
  assign \new_Sorter100|4173_  = \new_Sorter100|4073_  & \new_Sorter100|4074_ ;
  assign \new_Sorter100|4174_  = \new_Sorter100|4073_  | \new_Sorter100|4074_ ;
  assign \new_Sorter100|4175_  = \new_Sorter100|4075_  & \new_Sorter100|4076_ ;
  assign \new_Sorter100|4176_  = \new_Sorter100|4075_  | \new_Sorter100|4076_ ;
  assign \new_Sorter100|4177_  = \new_Sorter100|4077_  & \new_Sorter100|4078_ ;
  assign \new_Sorter100|4178_  = \new_Sorter100|4077_  | \new_Sorter100|4078_ ;
  assign \new_Sorter100|4179_  = \new_Sorter100|4079_  & \new_Sorter100|4080_ ;
  assign \new_Sorter100|4180_  = \new_Sorter100|4079_  | \new_Sorter100|4080_ ;
  assign \new_Sorter100|4181_  = \new_Sorter100|4081_  & \new_Sorter100|4082_ ;
  assign \new_Sorter100|4182_  = \new_Sorter100|4081_  | \new_Sorter100|4082_ ;
  assign \new_Sorter100|4183_  = \new_Sorter100|4083_  & \new_Sorter100|4084_ ;
  assign \new_Sorter100|4184_  = \new_Sorter100|4083_  | \new_Sorter100|4084_ ;
  assign \new_Sorter100|4185_  = \new_Sorter100|4085_  & \new_Sorter100|4086_ ;
  assign \new_Sorter100|4186_  = \new_Sorter100|4085_  | \new_Sorter100|4086_ ;
  assign \new_Sorter100|4187_  = \new_Sorter100|4087_  & \new_Sorter100|4088_ ;
  assign \new_Sorter100|4188_  = \new_Sorter100|4087_  | \new_Sorter100|4088_ ;
  assign \new_Sorter100|4189_  = \new_Sorter100|4089_  & \new_Sorter100|4090_ ;
  assign \new_Sorter100|4190_  = \new_Sorter100|4089_  | \new_Sorter100|4090_ ;
  assign \new_Sorter100|4191_  = \new_Sorter100|4091_  & \new_Sorter100|4092_ ;
  assign \new_Sorter100|4192_  = \new_Sorter100|4091_  | \new_Sorter100|4092_ ;
  assign \new_Sorter100|4193_  = \new_Sorter100|4093_  & \new_Sorter100|4094_ ;
  assign \new_Sorter100|4194_  = \new_Sorter100|4093_  | \new_Sorter100|4094_ ;
  assign \new_Sorter100|4195_  = \new_Sorter100|4095_  & \new_Sorter100|4096_ ;
  assign \new_Sorter100|4196_  = \new_Sorter100|4095_  | \new_Sorter100|4096_ ;
  assign \new_Sorter100|4197_  = \new_Sorter100|4097_  & \new_Sorter100|4098_ ;
  assign \new_Sorter100|4198_  = \new_Sorter100|4097_  | \new_Sorter100|4098_ ;
  assign \new_Sorter100|4200_  = \new_Sorter100|4100_  & \new_Sorter100|4101_ ;
  assign \new_Sorter100|4201_  = \new_Sorter100|4100_  | \new_Sorter100|4101_ ;
  assign \new_Sorter100|4202_  = \new_Sorter100|4102_  & \new_Sorter100|4103_ ;
  assign \new_Sorter100|4203_  = \new_Sorter100|4102_  | \new_Sorter100|4103_ ;
  assign \new_Sorter100|4204_  = \new_Sorter100|4104_  & \new_Sorter100|4105_ ;
  assign \new_Sorter100|4205_  = \new_Sorter100|4104_  | \new_Sorter100|4105_ ;
  assign \new_Sorter100|4206_  = \new_Sorter100|4106_  & \new_Sorter100|4107_ ;
  assign \new_Sorter100|4207_  = \new_Sorter100|4106_  | \new_Sorter100|4107_ ;
  assign \new_Sorter100|4208_  = \new_Sorter100|4108_  & \new_Sorter100|4109_ ;
  assign \new_Sorter100|4209_  = \new_Sorter100|4108_  | \new_Sorter100|4109_ ;
  assign \new_Sorter100|4210_  = \new_Sorter100|4110_  & \new_Sorter100|4111_ ;
  assign \new_Sorter100|4211_  = \new_Sorter100|4110_  | \new_Sorter100|4111_ ;
  assign \new_Sorter100|4212_  = \new_Sorter100|4112_  & \new_Sorter100|4113_ ;
  assign \new_Sorter100|4213_  = \new_Sorter100|4112_  | \new_Sorter100|4113_ ;
  assign \new_Sorter100|4214_  = \new_Sorter100|4114_  & \new_Sorter100|4115_ ;
  assign \new_Sorter100|4215_  = \new_Sorter100|4114_  | \new_Sorter100|4115_ ;
  assign \new_Sorter100|4216_  = \new_Sorter100|4116_  & \new_Sorter100|4117_ ;
  assign \new_Sorter100|4217_  = \new_Sorter100|4116_  | \new_Sorter100|4117_ ;
  assign \new_Sorter100|4218_  = \new_Sorter100|4118_  & \new_Sorter100|4119_ ;
  assign \new_Sorter100|4219_  = \new_Sorter100|4118_  | \new_Sorter100|4119_ ;
  assign \new_Sorter100|4220_  = \new_Sorter100|4120_  & \new_Sorter100|4121_ ;
  assign \new_Sorter100|4221_  = \new_Sorter100|4120_  | \new_Sorter100|4121_ ;
  assign \new_Sorter100|4222_  = \new_Sorter100|4122_  & \new_Sorter100|4123_ ;
  assign \new_Sorter100|4223_  = \new_Sorter100|4122_  | \new_Sorter100|4123_ ;
  assign \new_Sorter100|4224_  = \new_Sorter100|4124_  & \new_Sorter100|4125_ ;
  assign \new_Sorter100|4225_  = \new_Sorter100|4124_  | \new_Sorter100|4125_ ;
  assign \new_Sorter100|4226_  = \new_Sorter100|4126_  & \new_Sorter100|4127_ ;
  assign \new_Sorter100|4227_  = \new_Sorter100|4126_  | \new_Sorter100|4127_ ;
  assign \new_Sorter100|4228_  = \new_Sorter100|4128_  & \new_Sorter100|4129_ ;
  assign \new_Sorter100|4229_  = \new_Sorter100|4128_  | \new_Sorter100|4129_ ;
  assign \new_Sorter100|4230_  = \new_Sorter100|4130_  & \new_Sorter100|4131_ ;
  assign \new_Sorter100|4231_  = \new_Sorter100|4130_  | \new_Sorter100|4131_ ;
  assign \new_Sorter100|4232_  = \new_Sorter100|4132_  & \new_Sorter100|4133_ ;
  assign \new_Sorter100|4233_  = \new_Sorter100|4132_  | \new_Sorter100|4133_ ;
  assign \new_Sorter100|4234_  = \new_Sorter100|4134_  & \new_Sorter100|4135_ ;
  assign \new_Sorter100|4235_  = \new_Sorter100|4134_  | \new_Sorter100|4135_ ;
  assign \new_Sorter100|4236_  = \new_Sorter100|4136_  & \new_Sorter100|4137_ ;
  assign \new_Sorter100|4237_  = \new_Sorter100|4136_  | \new_Sorter100|4137_ ;
  assign \new_Sorter100|4238_  = \new_Sorter100|4138_  & \new_Sorter100|4139_ ;
  assign \new_Sorter100|4239_  = \new_Sorter100|4138_  | \new_Sorter100|4139_ ;
  assign \new_Sorter100|4240_  = \new_Sorter100|4140_  & \new_Sorter100|4141_ ;
  assign \new_Sorter100|4241_  = \new_Sorter100|4140_  | \new_Sorter100|4141_ ;
  assign \new_Sorter100|4242_  = \new_Sorter100|4142_  & \new_Sorter100|4143_ ;
  assign \new_Sorter100|4243_  = \new_Sorter100|4142_  | \new_Sorter100|4143_ ;
  assign \new_Sorter100|4244_  = \new_Sorter100|4144_  & \new_Sorter100|4145_ ;
  assign \new_Sorter100|4245_  = \new_Sorter100|4144_  | \new_Sorter100|4145_ ;
  assign \new_Sorter100|4246_  = \new_Sorter100|4146_  & \new_Sorter100|4147_ ;
  assign \new_Sorter100|4247_  = \new_Sorter100|4146_  | \new_Sorter100|4147_ ;
  assign \new_Sorter100|4248_  = \new_Sorter100|4148_  & \new_Sorter100|4149_ ;
  assign \new_Sorter100|4249_  = \new_Sorter100|4148_  | \new_Sorter100|4149_ ;
  assign \new_Sorter100|4250_  = \new_Sorter100|4150_  & \new_Sorter100|4151_ ;
  assign \new_Sorter100|4251_  = \new_Sorter100|4150_  | \new_Sorter100|4151_ ;
  assign \new_Sorter100|4252_  = \new_Sorter100|4152_  & \new_Sorter100|4153_ ;
  assign \new_Sorter100|4253_  = \new_Sorter100|4152_  | \new_Sorter100|4153_ ;
  assign \new_Sorter100|4254_  = \new_Sorter100|4154_  & \new_Sorter100|4155_ ;
  assign \new_Sorter100|4255_  = \new_Sorter100|4154_  | \new_Sorter100|4155_ ;
  assign \new_Sorter100|4256_  = \new_Sorter100|4156_  & \new_Sorter100|4157_ ;
  assign \new_Sorter100|4257_  = \new_Sorter100|4156_  | \new_Sorter100|4157_ ;
  assign \new_Sorter100|4258_  = \new_Sorter100|4158_  & \new_Sorter100|4159_ ;
  assign \new_Sorter100|4259_  = \new_Sorter100|4158_  | \new_Sorter100|4159_ ;
  assign \new_Sorter100|4260_  = \new_Sorter100|4160_  & \new_Sorter100|4161_ ;
  assign \new_Sorter100|4261_  = \new_Sorter100|4160_  | \new_Sorter100|4161_ ;
  assign \new_Sorter100|4262_  = \new_Sorter100|4162_  & \new_Sorter100|4163_ ;
  assign \new_Sorter100|4263_  = \new_Sorter100|4162_  | \new_Sorter100|4163_ ;
  assign \new_Sorter100|4264_  = \new_Sorter100|4164_  & \new_Sorter100|4165_ ;
  assign \new_Sorter100|4265_  = \new_Sorter100|4164_  | \new_Sorter100|4165_ ;
  assign \new_Sorter100|4266_  = \new_Sorter100|4166_  & \new_Sorter100|4167_ ;
  assign \new_Sorter100|4267_  = \new_Sorter100|4166_  | \new_Sorter100|4167_ ;
  assign \new_Sorter100|4268_  = \new_Sorter100|4168_  & \new_Sorter100|4169_ ;
  assign \new_Sorter100|4269_  = \new_Sorter100|4168_  | \new_Sorter100|4169_ ;
  assign \new_Sorter100|4270_  = \new_Sorter100|4170_  & \new_Sorter100|4171_ ;
  assign \new_Sorter100|4271_  = \new_Sorter100|4170_  | \new_Sorter100|4171_ ;
  assign \new_Sorter100|4272_  = \new_Sorter100|4172_  & \new_Sorter100|4173_ ;
  assign \new_Sorter100|4273_  = \new_Sorter100|4172_  | \new_Sorter100|4173_ ;
  assign \new_Sorter100|4274_  = \new_Sorter100|4174_  & \new_Sorter100|4175_ ;
  assign \new_Sorter100|4275_  = \new_Sorter100|4174_  | \new_Sorter100|4175_ ;
  assign \new_Sorter100|4276_  = \new_Sorter100|4176_  & \new_Sorter100|4177_ ;
  assign \new_Sorter100|4277_  = \new_Sorter100|4176_  | \new_Sorter100|4177_ ;
  assign \new_Sorter100|4278_  = \new_Sorter100|4178_  & \new_Sorter100|4179_ ;
  assign \new_Sorter100|4279_  = \new_Sorter100|4178_  | \new_Sorter100|4179_ ;
  assign \new_Sorter100|4280_  = \new_Sorter100|4180_  & \new_Sorter100|4181_ ;
  assign \new_Sorter100|4281_  = \new_Sorter100|4180_  | \new_Sorter100|4181_ ;
  assign \new_Sorter100|4282_  = \new_Sorter100|4182_  & \new_Sorter100|4183_ ;
  assign \new_Sorter100|4283_  = \new_Sorter100|4182_  | \new_Sorter100|4183_ ;
  assign \new_Sorter100|4284_  = \new_Sorter100|4184_  & \new_Sorter100|4185_ ;
  assign \new_Sorter100|4285_  = \new_Sorter100|4184_  | \new_Sorter100|4185_ ;
  assign \new_Sorter100|4286_  = \new_Sorter100|4186_  & \new_Sorter100|4187_ ;
  assign \new_Sorter100|4287_  = \new_Sorter100|4186_  | \new_Sorter100|4187_ ;
  assign \new_Sorter100|4288_  = \new_Sorter100|4188_  & \new_Sorter100|4189_ ;
  assign \new_Sorter100|4289_  = \new_Sorter100|4188_  | \new_Sorter100|4189_ ;
  assign \new_Sorter100|4290_  = \new_Sorter100|4190_  & \new_Sorter100|4191_ ;
  assign \new_Sorter100|4291_  = \new_Sorter100|4190_  | \new_Sorter100|4191_ ;
  assign \new_Sorter100|4292_  = \new_Sorter100|4192_  & \new_Sorter100|4193_ ;
  assign \new_Sorter100|4293_  = \new_Sorter100|4192_  | \new_Sorter100|4193_ ;
  assign \new_Sorter100|4294_  = \new_Sorter100|4194_  & \new_Sorter100|4195_ ;
  assign \new_Sorter100|4295_  = \new_Sorter100|4194_  | \new_Sorter100|4195_ ;
  assign \new_Sorter100|4296_  = \new_Sorter100|4196_  & \new_Sorter100|4197_ ;
  assign \new_Sorter100|4297_  = \new_Sorter100|4196_  | \new_Sorter100|4197_ ;
  assign \new_Sorter100|4298_  = \new_Sorter100|4198_  & \new_Sorter100|4199_ ;
  assign \new_Sorter100|4299_  = \new_Sorter100|4198_  | \new_Sorter100|4199_ ;
  assign \new_Sorter100|4300_  = \new_Sorter100|4200_ ;
  assign \new_Sorter100|4399_  = \new_Sorter100|4299_ ;
  assign \new_Sorter100|4301_  = \new_Sorter100|4201_  & \new_Sorter100|4202_ ;
  assign \new_Sorter100|4302_  = \new_Sorter100|4201_  | \new_Sorter100|4202_ ;
  assign \new_Sorter100|4303_  = \new_Sorter100|4203_  & \new_Sorter100|4204_ ;
  assign \new_Sorter100|4304_  = \new_Sorter100|4203_  | \new_Sorter100|4204_ ;
  assign \new_Sorter100|4305_  = \new_Sorter100|4205_  & \new_Sorter100|4206_ ;
  assign \new_Sorter100|4306_  = \new_Sorter100|4205_  | \new_Sorter100|4206_ ;
  assign \new_Sorter100|4307_  = \new_Sorter100|4207_  & \new_Sorter100|4208_ ;
  assign \new_Sorter100|4308_  = \new_Sorter100|4207_  | \new_Sorter100|4208_ ;
  assign \new_Sorter100|4309_  = \new_Sorter100|4209_  & \new_Sorter100|4210_ ;
  assign \new_Sorter100|4310_  = \new_Sorter100|4209_  | \new_Sorter100|4210_ ;
  assign \new_Sorter100|4311_  = \new_Sorter100|4211_  & \new_Sorter100|4212_ ;
  assign \new_Sorter100|4312_  = \new_Sorter100|4211_  | \new_Sorter100|4212_ ;
  assign \new_Sorter100|4313_  = \new_Sorter100|4213_  & \new_Sorter100|4214_ ;
  assign \new_Sorter100|4314_  = \new_Sorter100|4213_  | \new_Sorter100|4214_ ;
  assign \new_Sorter100|4315_  = \new_Sorter100|4215_  & \new_Sorter100|4216_ ;
  assign \new_Sorter100|4316_  = \new_Sorter100|4215_  | \new_Sorter100|4216_ ;
  assign \new_Sorter100|4317_  = \new_Sorter100|4217_  & \new_Sorter100|4218_ ;
  assign \new_Sorter100|4318_  = \new_Sorter100|4217_  | \new_Sorter100|4218_ ;
  assign \new_Sorter100|4319_  = \new_Sorter100|4219_  & \new_Sorter100|4220_ ;
  assign \new_Sorter100|4320_  = \new_Sorter100|4219_  | \new_Sorter100|4220_ ;
  assign \new_Sorter100|4321_  = \new_Sorter100|4221_  & \new_Sorter100|4222_ ;
  assign \new_Sorter100|4322_  = \new_Sorter100|4221_  | \new_Sorter100|4222_ ;
  assign \new_Sorter100|4323_  = \new_Sorter100|4223_  & \new_Sorter100|4224_ ;
  assign \new_Sorter100|4324_  = \new_Sorter100|4223_  | \new_Sorter100|4224_ ;
  assign \new_Sorter100|4325_  = \new_Sorter100|4225_  & \new_Sorter100|4226_ ;
  assign \new_Sorter100|4326_  = \new_Sorter100|4225_  | \new_Sorter100|4226_ ;
  assign \new_Sorter100|4327_  = \new_Sorter100|4227_  & \new_Sorter100|4228_ ;
  assign \new_Sorter100|4328_  = \new_Sorter100|4227_  | \new_Sorter100|4228_ ;
  assign \new_Sorter100|4329_  = \new_Sorter100|4229_  & \new_Sorter100|4230_ ;
  assign \new_Sorter100|4330_  = \new_Sorter100|4229_  | \new_Sorter100|4230_ ;
  assign \new_Sorter100|4331_  = \new_Sorter100|4231_  & \new_Sorter100|4232_ ;
  assign \new_Sorter100|4332_  = \new_Sorter100|4231_  | \new_Sorter100|4232_ ;
  assign \new_Sorter100|4333_  = \new_Sorter100|4233_  & \new_Sorter100|4234_ ;
  assign \new_Sorter100|4334_  = \new_Sorter100|4233_  | \new_Sorter100|4234_ ;
  assign \new_Sorter100|4335_  = \new_Sorter100|4235_  & \new_Sorter100|4236_ ;
  assign \new_Sorter100|4336_  = \new_Sorter100|4235_  | \new_Sorter100|4236_ ;
  assign \new_Sorter100|4337_  = \new_Sorter100|4237_  & \new_Sorter100|4238_ ;
  assign \new_Sorter100|4338_  = \new_Sorter100|4237_  | \new_Sorter100|4238_ ;
  assign \new_Sorter100|4339_  = \new_Sorter100|4239_  & \new_Sorter100|4240_ ;
  assign \new_Sorter100|4340_  = \new_Sorter100|4239_  | \new_Sorter100|4240_ ;
  assign \new_Sorter100|4341_  = \new_Sorter100|4241_  & \new_Sorter100|4242_ ;
  assign \new_Sorter100|4342_  = \new_Sorter100|4241_  | \new_Sorter100|4242_ ;
  assign \new_Sorter100|4343_  = \new_Sorter100|4243_  & \new_Sorter100|4244_ ;
  assign \new_Sorter100|4344_  = \new_Sorter100|4243_  | \new_Sorter100|4244_ ;
  assign \new_Sorter100|4345_  = \new_Sorter100|4245_  & \new_Sorter100|4246_ ;
  assign \new_Sorter100|4346_  = \new_Sorter100|4245_  | \new_Sorter100|4246_ ;
  assign \new_Sorter100|4347_  = \new_Sorter100|4247_  & \new_Sorter100|4248_ ;
  assign \new_Sorter100|4348_  = \new_Sorter100|4247_  | \new_Sorter100|4248_ ;
  assign \new_Sorter100|4349_  = \new_Sorter100|4249_  & \new_Sorter100|4250_ ;
  assign \new_Sorter100|4350_  = \new_Sorter100|4249_  | \new_Sorter100|4250_ ;
  assign \new_Sorter100|4351_  = \new_Sorter100|4251_  & \new_Sorter100|4252_ ;
  assign \new_Sorter100|4352_  = \new_Sorter100|4251_  | \new_Sorter100|4252_ ;
  assign \new_Sorter100|4353_  = \new_Sorter100|4253_  & \new_Sorter100|4254_ ;
  assign \new_Sorter100|4354_  = \new_Sorter100|4253_  | \new_Sorter100|4254_ ;
  assign \new_Sorter100|4355_  = \new_Sorter100|4255_  & \new_Sorter100|4256_ ;
  assign \new_Sorter100|4356_  = \new_Sorter100|4255_  | \new_Sorter100|4256_ ;
  assign \new_Sorter100|4357_  = \new_Sorter100|4257_  & \new_Sorter100|4258_ ;
  assign \new_Sorter100|4358_  = \new_Sorter100|4257_  | \new_Sorter100|4258_ ;
  assign \new_Sorter100|4359_  = \new_Sorter100|4259_  & \new_Sorter100|4260_ ;
  assign \new_Sorter100|4360_  = \new_Sorter100|4259_  | \new_Sorter100|4260_ ;
  assign \new_Sorter100|4361_  = \new_Sorter100|4261_  & \new_Sorter100|4262_ ;
  assign \new_Sorter100|4362_  = \new_Sorter100|4261_  | \new_Sorter100|4262_ ;
  assign \new_Sorter100|4363_  = \new_Sorter100|4263_  & \new_Sorter100|4264_ ;
  assign \new_Sorter100|4364_  = \new_Sorter100|4263_  | \new_Sorter100|4264_ ;
  assign \new_Sorter100|4365_  = \new_Sorter100|4265_  & \new_Sorter100|4266_ ;
  assign \new_Sorter100|4366_  = \new_Sorter100|4265_  | \new_Sorter100|4266_ ;
  assign \new_Sorter100|4367_  = \new_Sorter100|4267_  & \new_Sorter100|4268_ ;
  assign \new_Sorter100|4368_  = \new_Sorter100|4267_  | \new_Sorter100|4268_ ;
  assign \new_Sorter100|4369_  = \new_Sorter100|4269_  & \new_Sorter100|4270_ ;
  assign \new_Sorter100|4370_  = \new_Sorter100|4269_  | \new_Sorter100|4270_ ;
  assign \new_Sorter100|4371_  = \new_Sorter100|4271_  & \new_Sorter100|4272_ ;
  assign \new_Sorter100|4372_  = \new_Sorter100|4271_  | \new_Sorter100|4272_ ;
  assign \new_Sorter100|4373_  = \new_Sorter100|4273_  & \new_Sorter100|4274_ ;
  assign \new_Sorter100|4374_  = \new_Sorter100|4273_  | \new_Sorter100|4274_ ;
  assign \new_Sorter100|4375_  = \new_Sorter100|4275_  & \new_Sorter100|4276_ ;
  assign \new_Sorter100|4376_  = \new_Sorter100|4275_  | \new_Sorter100|4276_ ;
  assign \new_Sorter100|4377_  = \new_Sorter100|4277_  & \new_Sorter100|4278_ ;
  assign \new_Sorter100|4378_  = \new_Sorter100|4277_  | \new_Sorter100|4278_ ;
  assign \new_Sorter100|4379_  = \new_Sorter100|4279_  & \new_Sorter100|4280_ ;
  assign \new_Sorter100|4380_  = \new_Sorter100|4279_  | \new_Sorter100|4280_ ;
  assign \new_Sorter100|4381_  = \new_Sorter100|4281_  & \new_Sorter100|4282_ ;
  assign \new_Sorter100|4382_  = \new_Sorter100|4281_  | \new_Sorter100|4282_ ;
  assign \new_Sorter100|4383_  = \new_Sorter100|4283_  & \new_Sorter100|4284_ ;
  assign \new_Sorter100|4384_  = \new_Sorter100|4283_  | \new_Sorter100|4284_ ;
  assign \new_Sorter100|4385_  = \new_Sorter100|4285_  & \new_Sorter100|4286_ ;
  assign \new_Sorter100|4386_  = \new_Sorter100|4285_  | \new_Sorter100|4286_ ;
  assign \new_Sorter100|4387_  = \new_Sorter100|4287_  & \new_Sorter100|4288_ ;
  assign \new_Sorter100|4388_  = \new_Sorter100|4287_  | \new_Sorter100|4288_ ;
  assign \new_Sorter100|4389_  = \new_Sorter100|4289_  & \new_Sorter100|4290_ ;
  assign \new_Sorter100|4390_  = \new_Sorter100|4289_  | \new_Sorter100|4290_ ;
  assign \new_Sorter100|4391_  = \new_Sorter100|4291_  & \new_Sorter100|4292_ ;
  assign \new_Sorter100|4392_  = \new_Sorter100|4291_  | \new_Sorter100|4292_ ;
  assign \new_Sorter100|4393_  = \new_Sorter100|4293_  & \new_Sorter100|4294_ ;
  assign \new_Sorter100|4394_  = \new_Sorter100|4293_  | \new_Sorter100|4294_ ;
  assign \new_Sorter100|4395_  = \new_Sorter100|4295_  & \new_Sorter100|4296_ ;
  assign \new_Sorter100|4396_  = \new_Sorter100|4295_  | \new_Sorter100|4296_ ;
  assign \new_Sorter100|4397_  = \new_Sorter100|4297_  & \new_Sorter100|4298_ ;
  assign \new_Sorter100|4398_  = \new_Sorter100|4297_  | \new_Sorter100|4298_ ;
  assign \new_Sorter100|4400_  = \new_Sorter100|4300_  & \new_Sorter100|4301_ ;
  assign \new_Sorter100|4401_  = \new_Sorter100|4300_  | \new_Sorter100|4301_ ;
  assign \new_Sorter100|4402_  = \new_Sorter100|4302_  & \new_Sorter100|4303_ ;
  assign \new_Sorter100|4403_  = \new_Sorter100|4302_  | \new_Sorter100|4303_ ;
  assign \new_Sorter100|4404_  = \new_Sorter100|4304_  & \new_Sorter100|4305_ ;
  assign \new_Sorter100|4405_  = \new_Sorter100|4304_  | \new_Sorter100|4305_ ;
  assign \new_Sorter100|4406_  = \new_Sorter100|4306_  & \new_Sorter100|4307_ ;
  assign \new_Sorter100|4407_  = \new_Sorter100|4306_  | \new_Sorter100|4307_ ;
  assign \new_Sorter100|4408_  = \new_Sorter100|4308_  & \new_Sorter100|4309_ ;
  assign \new_Sorter100|4409_  = \new_Sorter100|4308_  | \new_Sorter100|4309_ ;
  assign \new_Sorter100|4410_  = \new_Sorter100|4310_  & \new_Sorter100|4311_ ;
  assign \new_Sorter100|4411_  = \new_Sorter100|4310_  | \new_Sorter100|4311_ ;
  assign \new_Sorter100|4412_  = \new_Sorter100|4312_  & \new_Sorter100|4313_ ;
  assign \new_Sorter100|4413_  = \new_Sorter100|4312_  | \new_Sorter100|4313_ ;
  assign \new_Sorter100|4414_  = \new_Sorter100|4314_  & \new_Sorter100|4315_ ;
  assign \new_Sorter100|4415_  = \new_Sorter100|4314_  | \new_Sorter100|4315_ ;
  assign \new_Sorter100|4416_  = \new_Sorter100|4316_  & \new_Sorter100|4317_ ;
  assign \new_Sorter100|4417_  = \new_Sorter100|4316_  | \new_Sorter100|4317_ ;
  assign \new_Sorter100|4418_  = \new_Sorter100|4318_  & \new_Sorter100|4319_ ;
  assign \new_Sorter100|4419_  = \new_Sorter100|4318_  | \new_Sorter100|4319_ ;
  assign \new_Sorter100|4420_  = \new_Sorter100|4320_  & \new_Sorter100|4321_ ;
  assign \new_Sorter100|4421_  = \new_Sorter100|4320_  | \new_Sorter100|4321_ ;
  assign \new_Sorter100|4422_  = \new_Sorter100|4322_  & \new_Sorter100|4323_ ;
  assign \new_Sorter100|4423_  = \new_Sorter100|4322_  | \new_Sorter100|4323_ ;
  assign \new_Sorter100|4424_  = \new_Sorter100|4324_  & \new_Sorter100|4325_ ;
  assign \new_Sorter100|4425_  = \new_Sorter100|4324_  | \new_Sorter100|4325_ ;
  assign \new_Sorter100|4426_  = \new_Sorter100|4326_  & \new_Sorter100|4327_ ;
  assign \new_Sorter100|4427_  = \new_Sorter100|4326_  | \new_Sorter100|4327_ ;
  assign \new_Sorter100|4428_  = \new_Sorter100|4328_  & \new_Sorter100|4329_ ;
  assign \new_Sorter100|4429_  = \new_Sorter100|4328_  | \new_Sorter100|4329_ ;
  assign \new_Sorter100|4430_  = \new_Sorter100|4330_  & \new_Sorter100|4331_ ;
  assign \new_Sorter100|4431_  = \new_Sorter100|4330_  | \new_Sorter100|4331_ ;
  assign \new_Sorter100|4432_  = \new_Sorter100|4332_  & \new_Sorter100|4333_ ;
  assign \new_Sorter100|4433_  = \new_Sorter100|4332_  | \new_Sorter100|4333_ ;
  assign \new_Sorter100|4434_  = \new_Sorter100|4334_  & \new_Sorter100|4335_ ;
  assign \new_Sorter100|4435_  = \new_Sorter100|4334_  | \new_Sorter100|4335_ ;
  assign \new_Sorter100|4436_  = \new_Sorter100|4336_  & \new_Sorter100|4337_ ;
  assign \new_Sorter100|4437_  = \new_Sorter100|4336_  | \new_Sorter100|4337_ ;
  assign \new_Sorter100|4438_  = \new_Sorter100|4338_  & \new_Sorter100|4339_ ;
  assign \new_Sorter100|4439_  = \new_Sorter100|4338_  | \new_Sorter100|4339_ ;
  assign \new_Sorter100|4440_  = \new_Sorter100|4340_  & \new_Sorter100|4341_ ;
  assign \new_Sorter100|4441_  = \new_Sorter100|4340_  | \new_Sorter100|4341_ ;
  assign \new_Sorter100|4442_  = \new_Sorter100|4342_  & \new_Sorter100|4343_ ;
  assign \new_Sorter100|4443_  = \new_Sorter100|4342_  | \new_Sorter100|4343_ ;
  assign \new_Sorter100|4444_  = \new_Sorter100|4344_  & \new_Sorter100|4345_ ;
  assign \new_Sorter100|4445_  = \new_Sorter100|4344_  | \new_Sorter100|4345_ ;
  assign \new_Sorter100|4446_  = \new_Sorter100|4346_  & \new_Sorter100|4347_ ;
  assign \new_Sorter100|4447_  = \new_Sorter100|4346_  | \new_Sorter100|4347_ ;
  assign \new_Sorter100|4448_  = \new_Sorter100|4348_  & \new_Sorter100|4349_ ;
  assign \new_Sorter100|4449_  = \new_Sorter100|4348_  | \new_Sorter100|4349_ ;
  assign \new_Sorter100|4450_  = \new_Sorter100|4350_  & \new_Sorter100|4351_ ;
  assign \new_Sorter100|4451_  = \new_Sorter100|4350_  | \new_Sorter100|4351_ ;
  assign \new_Sorter100|4452_  = \new_Sorter100|4352_  & \new_Sorter100|4353_ ;
  assign \new_Sorter100|4453_  = \new_Sorter100|4352_  | \new_Sorter100|4353_ ;
  assign \new_Sorter100|4454_  = \new_Sorter100|4354_  & \new_Sorter100|4355_ ;
  assign \new_Sorter100|4455_  = \new_Sorter100|4354_  | \new_Sorter100|4355_ ;
  assign \new_Sorter100|4456_  = \new_Sorter100|4356_  & \new_Sorter100|4357_ ;
  assign \new_Sorter100|4457_  = \new_Sorter100|4356_  | \new_Sorter100|4357_ ;
  assign \new_Sorter100|4458_  = \new_Sorter100|4358_  & \new_Sorter100|4359_ ;
  assign \new_Sorter100|4459_  = \new_Sorter100|4358_  | \new_Sorter100|4359_ ;
  assign \new_Sorter100|4460_  = \new_Sorter100|4360_  & \new_Sorter100|4361_ ;
  assign \new_Sorter100|4461_  = \new_Sorter100|4360_  | \new_Sorter100|4361_ ;
  assign \new_Sorter100|4462_  = \new_Sorter100|4362_  & \new_Sorter100|4363_ ;
  assign \new_Sorter100|4463_  = \new_Sorter100|4362_  | \new_Sorter100|4363_ ;
  assign \new_Sorter100|4464_  = \new_Sorter100|4364_  & \new_Sorter100|4365_ ;
  assign \new_Sorter100|4465_  = \new_Sorter100|4364_  | \new_Sorter100|4365_ ;
  assign \new_Sorter100|4466_  = \new_Sorter100|4366_  & \new_Sorter100|4367_ ;
  assign \new_Sorter100|4467_  = \new_Sorter100|4366_  | \new_Sorter100|4367_ ;
  assign \new_Sorter100|4468_  = \new_Sorter100|4368_  & \new_Sorter100|4369_ ;
  assign \new_Sorter100|4469_  = \new_Sorter100|4368_  | \new_Sorter100|4369_ ;
  assign \new_Sorter100|4470_  = \new_Sorter100|4370_  & \new_Sorter100|4371_ ;
  assign \new_Sorter100|4471_  = \new_Sorter100|4370_  | \new_Sorter100|4371_ ;
  assign \new_Sorter100|4472_  = \new_Sorter100|4372_  & \new_Sorter100|4373_ ;
  assign \new_Sorter100|4473_  = \new_Sorter100|4372_  | \new_Sorter100|4373_ ;
  assign \new_Sorter100|4474_  = \new_Sorter100|4374_  & \new_Sorter100|4375_ ;
  assign \new_Sorter100|4475_  = \new_Sorter100|4374_  | \new_Sorter100|4375_ ;
  assign \new_Sorter100|4476_  = \new_Sorter100|4376_  & \new_Sorter100|4377_ ;
  assign \new_Sorter100|4477_  = \new_Sorter100|4376_  | \new_Sorter100|4377_ ;
  assign \new_Sorter100|4478_  = \new_Sorter100|4378_  & \new_Sorter100|4379_ ;
  assign \new_Sorter100|4479_  = \new_Sorter100|4378_  | \new_Sorter100|4379_ ;
  assign \new_Sorter100|4480_  = \new_Sorter100|4380_  & \new_Sorter100|4381_ ;
  assign \new_Sorter100|4481_  = \new_Sorter100|4380_  | \new_Sorter100|4381_ ;
  assign \new_Sorter100|4482_  = \new_Sorter100|4382_  & \new_Sorter100|4383_ ;
  assign \new_Sorter100|4483_  = \new_Sorter100|4382_  | \new_Sorter100|4383_ ;
  assign \new_Sorter100|4484_  = \new_Sorter100|4384_  & \new_Sorter100|4385_ ;
  assign \new_Sorter100|4485_  = \new_Sorter100|4384_  | \new_Sorter100|4385_ ;
  assign \new_Sorter100|4486_  = \new_Sorter100|4386_  & \new_Sorter100|4387_ ;
  assign \new_Sorter100|4487_  = \new_Sorter100|4386_  | \new_Sorter100|4387_ ;
  assign \new_Sorter100|4488_  = \new_Sorter100|4388_  & \new_Sorter100|4389_ ;
  assign \new_Sorter100|4489_  = \new_Sorter100|4388_  | \new_Sorter100|4389_ ;
  assign \new_Sorter100|4490_  = \new_Sorter100|4390_  & \new_Sorter100|4391_ ;
  assign \new_Sorter100|4491_  = \new_Sorter100|4390_  | \new_Sorter100|4391_ ;
  assign \new_Sorter100|4492_  = \new_Sorter100|4392_  & \new_Sorter100|4393_ ;
  assign \new_Sorter100|4493_  = \new_Sorter100|4392_  | \new_Sorter100|4393_ ;
  assign \new_Sorter100|4494_  = \new_Sorter100|4394_  & \new_Sorter100|4395_ ;
  assign \new_Sorter100|4495_  = \new_Sorter100|4394_  | \new_Sorter100|4395_ ;
  assign \new_Sorter100|4496_  = \new_Sorter100|4396_  & \new_Sorter100|4397_ ;
  assign \new_Sorter100|4497_  = \new_Sorter100|4396_  | \new_Sorter100|4397_ ;
  assign \new_Sorter100|4498_  = \new_Sorter100|4398_  & \new_Sorter100|4399_ ;
  assign \new_Sorter100|4499_  = \new_Sorter100|4398_  | \new_Sorter100|4399_ ;
  assign \new_Sorter100|4500_  = \new_Sorter100|4400_ ;
  assign \new_Sorter100|4599_  = \new_Sorter100|4499_ ;
  assign \new_Sorter100|4501_  = \new_Sorter100|4401_  & \new_Sorter100|4402_ ;
  assign \new_Sorter100|4502_  = \new_Sorter100|4401_  | \new_Sorter100|4402_ ;
  assign \new_Sorter100|4503_  = \new_Sorter100|4403_  & \new_Sorter100|4404_ ;
  assign \new_Sorter100|4504_  = \new_Sorter100|4403_  | \new_Sorter100|4404_ ;
  assign \new_Sorter100|4505_  = \new_Sorter100|4405_  & \new_Sorter100|4406_ ;
  assign \new_Sorter100|4506_  = \new_Sorter100|4405_  | \new_Sorter100|4406_ ;
  assign \new_Sorter100|4507_  = \new_Sorter100|4407_  & \new_Sorter100|4408_ ;
  assign \new_Sorter100|4508_  = \new_Sorter100|4407_  | \new_Sorter100|4408_ ;
  assign \new_Sorter100|4509_  = \new_Sorter100|4409_  & \new_Sorter100|4410_ ;
  assign \new_Sorter100|4510_  = \new_Sorter100|4409_  | \new_Sorter100|4410_ ;
  assign \new_Sorter100|4511_  = \new_Sorter100|4411_  & \new_Sorter100|4412_ ;
  assign \new_Sorter100|4512_  = \new_Sorter100|4411_  | \new_Sorter100|4412_ ;
  assign \new_Sorter100|4513_  = \new_Sorter100|4413_  & \new_Sorter100|4414_ ;
  assign \new_Sorter100|4514_  = \new_Sorter100|4413_  | \new_Sorter100|4414_ ;
  assign \new_Sorter100|4515_  = \new_Sorter100|4415_  & \new_Sorter100|4416_ ;
  assign \new_Sorter100|4516_  = \new_Sorter100|4415_  | \new_Sorter100|4416_ ;
  assign \new_Sorter100|4517_  = \new_Sorter100|4417_  & \new_Sorter100|4418_ ;
  assign \new_Sorter100|4518_  = \new_Sorter100|4417_  | \new_Sorter100|4418_ ;
  assign \new_Sorter100|4519_  = \new_Sorter100|4419_  & \new_Sorter100|4420_ ;
  assign \new_Sorter100|4520_  = \new_Sorter100|4419_  | \new_Sorter100|4420_ ;
  assign \new_Sorter100|4521_  = \new_Sorter100|4421_  & \new_Sorter100|4422_ ;
  assign \new_Sorter100|4522_  = \new_Sorter100|4421_  | \new_Sorter100|4422_ ;
  assign \new_Sorter100|4523_  = \new_Sorter100|4423_  & \new_Sorter100|4424_ ;
  assign \new_Sorter100|4524_  = \new_Sorter100|4423_  | \new_Sorter100|4424_ ;
  assign \new_Sorter100|4525_  = \new_Sorter100|4425_  & \new_Sorter100|4426_ ;
  assign \new_Sorter100|4526_  = \new_Sorter100|4425_  | \new_Sorter100|4426_ ;
  assign \new_Sorter100|4527_  = \new_Sorter100|4427_  & \new_Sorter100|4428_ ;
  assign \new_Sorter100|4528_  = \new_Sorter100|4427_  | \new_Sorter100|4428_ ;
  assign \new_Sorter100|4529_  = \new_Sorter100|4429_  & \new_Sorter100|4430_ ;
  assign \new_Sorter100|4530_  = \new_Sorter100|4429_  | \new_Sorter100|4430_ ;
  assign \new_Sorter100|4531_  = \new_Sorter100|4431_  & \new_Sorter100|4432_ ;
  assign \new_Sorter100|4532_  = \new_Sorter100|4431_  | \new_Sorter100|4432_ ;
  assign \new_Sorter100|4533_  = \new_Sorter100|4433_  & \new_Sorter100|4434_ ;
  assign \new_Sorter100|4534_  = \new_Sorter100|4433_  | \new_Sorter100|4434_ ;
  assign \new_Sorter100|4535_  = \new_Sorter100|4435_  & \new_Sorter100|4436_ ;
  assign \new_Sorter100|4536_  = \new_Sorter100|4435_  | \new_Sorter100|4436_ ;
  assign \new_Sorter100|4537_  = \new_Sorter100|4437_  & \new_Sorter100|4438_ ;
  assign \new_Sorter100|4538_  = \new_Sorter100|4437_  | \new_Sorter100|4438_ ;
  assign \new_Sorter100|4539_  = \new_Sorter100|4439_  & \new_Sorter100|4440_ ;
  assign \new_Sorter100|4540_  = \new_Sorter100|4439_  | \new_Sorter100|4440_ ;
  assign \new_Sorter100|4541_  = \new_Sorter100|4441_  & \new_Sorter100|4442_ ;
  assign \new_Sorter100|4542_  = \new_Sorter100|4441_  | \new_Sorter100|4442_ ;
  assign \new_Sorter100|4543_  = \new_Sorter100|4443_  & \new_Sorter100|4444_ ;
  assign \new_Sorter100|4544_  = \new_Sorter100|4443_  | \new_Sorter100|4444_ ;
  assign \new_Sorter100|4545_  = \new_Sorter100|4445_  & \new_Sorter100|4446_ ;
  assign \new_Sorter100|4546_  = \new_Sorter100|4445_  | \new_Sorter100|4446_ ;
  assign \new_Sorter100|4547_  = \new_Sorter100|4447_  & \new_Sorter100|4448_ ;
  assign \new_Sorter100|4548_  = \new_Sorter100|4447_  | \new_Sorter100|4448_ ;
  assign \new_Sorter100|4549_  = \new_Sorter100|4449_  & \new_Sorter100|4450_ ;
  assign \new_Sorter100|4550_  = \new_Sorter100|4449_  | \new_Sorter100|4450_ ;
  assign \new_Sorter100|4551_  = \new_Sorter100|4451_  & \new_Sorter100|4452_ ;
  assign \new_Sorter100|4552_  = \new_Sorter100|4451_  | \new_Sorter100|4452_ ;
  assign \new_Sorter100|4553_  = \new_Sorter100|4453_  & \new_Sorter100|4454_ ;
  assign \new_Sorter100|4554_  = \new_Sorter100|4453_  | \new_Sorter100|4454_ ;
  assign \new_Sorter100|4555_  = \new_Sorter100|4455_  & \new_Sorter100|4456_ ;
  assign \new_Sorter100|4556_  = \new_Sorter100|4455_  | \new_Sorter100|4456_ ;
  assign \new_Sorter100|4557_  = \new_Sorter100|4457_  & \new_Sorter100|4458_ ;
  assign \new_Sorter100|4558_  = \new_Sorter100|4457_  | \new_Sorter100|4458_ ;
  assign \new_Sorter100|4559_  = \new_Sorter100|4459_  & \new_Sorter100|4460_ ;
  assign \new_Sorter100|4560_  = \new_Sorter100|4459_  | \new_Sorter100|4460_ ;
  assign \new_Sorter100|4561_  = \new_Sorter100|4461_  & \new_Sorter100|4462_ ;
  assign \new_Sorter100|4562_  = \new_Sorter100|4461_  | \new_Sorter100|4462_ ;
  assign \new_Sorter100|4563_  = \new_Sorter100|4463_  & \new_Sorter100|4464_ ;
  assign \new_Sorter100|4564_  = \new_Sorter100|4463_  | \new_Sorter100|4464_ ;
  assign \new_Sorter100|4565_  = \new_Sorter100|4465_  & \new_Sorter100|4466_ ;
  assign \new_Sorter100|4566_  = \new_Sorter100|4465_  | \new_Sorter100|4466_ ;
  assign \new_Sorter100|4567_  = \new_Sorter100|4467_  & \new_Sorter100|4468_ ;
  assign \new_Sorter100|4568_  = \new_Sorter100|4467_  | \new_Sorter100|4468_ ;
  assign \new_Sorter100|4569_  = \new_Sorter100|4469_  & \new_Sorter100|4470_ ;
  assign \new_Sorter100|4570_  = \new_Sorter100|4469_  | \new_Sorter100|4470_ ;
  assign \new_Sorter100|4571_  = \new_Sorter100|4471_  & \new_Sorter100|4472_ ;
  assign \new_Sorter100|4572_  = \new_Sorter100|4471_  | \new_Sorter100|4472_ ;
  assign \new_Sorter100|4573_  = \new_Sorter100|4473_  & \new_Sorter100|4474_ ;
  assign \new_Sorter100|4574_  = \new_Sorter100|4473_  | \new_Sorter100|4474_ ;
  assign \new_Sorter100|4575_  = \new_Sorter100|4475_  & \new_Sorter100|4476_ ;
  assign \new_Sorter100|4576_  = \new_Sorter100|4475_  | \new_Sorter100|4476_ ;
  assign \new_Sorter100|4577_  = \new_Sorter100|4477_  & \new_Sorter100|4478_ ;
  assign \new_Sorter100|4578_  = \new_Sorter100|4477_  | \new_Sorter100|4478_ ;
  assign \new_Sorter100|4579_  = \new_Sorter100|4479_  & \new_Sorter100|4480_ ;
  assign \new_Sorter100|4580_  = \new_Sorter100|4479_  | \new_Sorter100|4480_ ;
  assign \new_Sorter100|4581_  = \new_Sorter100|4481_  & \new_Sorter100|4482_ ;
  assign \new_Sorter100|4582_  = \new_Sorter100|4481_  | \new_Sorter100|4482_ ;
  assign \new_Sorter100|4583_  = \new_Sorter100|4483_  & \new_Sorter100|4484_ ;
  assign \new_Sorter100|4584_  = \new_Sorter100|4483_  | \new_Sorter100|4484_ ;
  assign \new_Sorter100|4585_  = \new_Sorter100|4485_  & \new_Sorter100|4486_ ;
  assign \new_Sorter100|4586_  = \new_Sorter100|4485_  | \new_Sorter100|4486_ ;
  assign \new_Sorter100|4587_  = \new_Sorter100|4487_  & \new_Sorter100|4488_ ;
  assign \new_Sorter100|4588_  = \new_Sorter100|4487_  | \new_Sorter100|4488_ ;
  assign \new_Sorter100|4589_  = \new_Sorter100|4489_  & \new_Sorter100|4490_ ;
  assign \new_Sorter100|4590_  = \new_Sorter100|4489_  | \new_Sorter100|4490_ ;
  assign \new_Sorter100|4591_  = \new_Sorter100|4491_  & \new_Sorter100|4492_ ;
  assign \new_Sorter100|4592_  = \new_Sorter100|4491_  | \new_Sorter100|4492_ ;
  assign \new_Sorter100|4593_  = \new_Sorter100|4493_  & \new_Sorter100|4494_ ;
  assign \new_Sorter100|4594_  = \new_Sorter100|4493_  | \new_Sorter100|4494_ ;
  assign \new_Sorter100|4595_  = \new_Sorter100|4495_  & \new_Sorter100|4496_ ;
  assign \new_Sorter100|4596_  = \new_Sorter100|4495_  | \new_Sorter100|4496_ ;
  assign \new_Sorter100|4597_  = \new_Sorter100|4497_  & \new_Sorter100|4498_ ;
  assign \new_Sorter100|4598_  = \new_Sorter100|4497_  | \new_Sorter100|4498_ ;
  assign \new_Sorter100|4600_  = \new_Sorter100|4500_  & \new_Sorter100|4501_ ;
  assign \new_Sorter100|4601_  = \new_Sorter100|4500_  | \new_Sorter100|4501_ ;
  assign \new_Sorter100|4602_  = \new_Sorter100|4502_  & \new_Sorter100|4503_ ;
  assign \new_Sorter100|4603_  = \new_Sorter100|4502_  | \new_Sorter100|4503_ ;
  assign \new_Sorter100|4604_  = \new_Sorter100|4504_  & \new_Sorter100|4505_ ;
  assign \new_Sorter100|4605_  = \new_Sorter100|4504_  | \new_Sorter100|4505_ ;
  assign \new_Sorter100|4606_  = \new_Sorter100|4506_  & \new_Sorter100|4507_ ;
  assign \new_Sorter100|4607_  = \new_Sorter100|4506_  | \new_Sorter100|4507_ ;
  assign \new_Sorter100|4608_  = \new_Sorter100|4508_  & \new_Sorter100|4509_ ;
  assign \new_Sorter100|4609_  = \new_Sorter100|4508_  | \new_Sorter100|4509_ ;
  assign \new_Sorter100|4610_  = \new_Sorter100|4510_  & \new_Sorter100|4511_ ;
  assign \new_Sorter100|4611_  = \new_Sorter100|4510_  | \new_Sorter100|4511_ ;
  assign \new_Sorter100|4612_  = \new_Sorter100|4512_  & \new_Sorter100|4513_ ;
  assign \new_Sorter100|4613_  = \new_Sorter100|4512_  | \new_Sorter100|4513_ ;
  assign \new_Sorter100|4614_  = \new_Sorter100|4514_  & \new_Sorter100|4515_ ;
  assign \new_Sorter100|4615_  = \new_Sorter100|4514_  | \new_Sorter100|4515_ ;
  assign \new_Sorter100|4616_  = \new_Sorter100|4516_  & \new_Sorter100|4517_ ;
  assign \new_Sorter100|4617_  = \new_Sorter100|4516_  | \new_Sorter100|4517_ ;
  assign \new_Sorter100|4618_  = \new_Sorter100|4518_  & \new_Sorter100|4519_ ;
  assign \new_Sorter100|4619_  = \new_Sorter100|4518_  | \new_Sorter100|4519_ ;
  assign \new_Sorter100|4620_  = \new_Sorter100|4520_  & \new_Sorter100|4521_ ;
  assign \new_Sorter100|4621_  = \new_Sorter100|4520_  | \new_Sorter100|4521_ ;
  assign \new_Sorter100|4622_  = \new_Sorter100|4522_  & \new_Sorter100|4523_ ;
  assign \new_Sorter100|4623_  = \new_Sorter100|4522_  | \new_Sorter100|4523_ ;
  assign \new_Sorter100|4624_  = \new_Sorter100|4524_  & \new_Sorter100|4525_ ;
  assign \new_Sorter100|4625_  = \new_Sorter100|4524_  | \new_Sorter100|4525_ ;
  assign \new_Sorter100|4626_  = \new_Sorter100|4526_  & \new_Sorter100|4527_ ;
  assign \new_Sorter100|4627_  = \new_Sorter100|4526_  | \new_Sorter100|4527_ ;
  assign \new_Sorter100|4628_  = \new_Sorter100|4528_  & \new_Sorter100|4529_ ;
  assign \new_Sorter100|4629_  = \new_Sorter100|4528_  | \new_Sorter100|4529_ ;
  assign \new_Sorter100|4630_  = \new_Sorter100|4530_  & \new_Sorter100|4531_ ;
  assign \new_Sorter100|4631_  = \new_Sorter100|4530_  | \new_Sorter100|4531_ ;
  assign \new_Sorter100|4632_  = \new_Sorter100|4532_  & \new_Sorter100|4533_ ;
  assign \new_Sorter100|4633_  = \new_Sorter100|4532_  | \new_Sorter100|4533_ ;
  assign \new_Sorter100|4634_  = \new_Sorter100|4534_  & \new_Sorter100|4535_ ;
  assign \new_Sorter100|4635_  = \new_Sorter100|4534_  | \new_Sorter100|4535_ ;
  assign \new_Sorter100|4636_  = \new_Sorter100|4536_  & \new_Sorter100|4537_ ;
  assign \new_Sorter100|4637_  = \new_Sorter100|4536_  | \new_Sorter100|4537_ ;
  assign \new_Sorter100|4638_  = \new_Sorter100|4538_  & \new_Sorter100|4539_ ;
  assign \new_Sorter100|4639_  = \new_Sorter100|4538_  | \new_Sorter100|4539_ ;
  assign \new_Sorter100|4640_  = \new_Sorter100|4540_  & \new_Sorter100|4541_ ;
  assign \new_Sorter100|4641_  = \new_Sorter100|4540_  | \new_Sorter100|4541_ ;
  assign \new_Sorter100|4642_  = \new_Sorter100|4542_  & \new_Sorter100|4543_ ;
  assign \new_Sorter100|4643_  = \new_Sorter100|4542_  | \new_Sorter100|4543_ ;
  assign \new_Sorter100|4644_  = \new_Sorter100|4544_  & \new_Sorter100|4545_ ;
  assign \new_Sorter100|4645_  = \new_Sorter100|4544_  | \new_Sorter100|4545_ ;
  assign \new_Sorter100|4646_  = \new_Sorter100|4546_  & \new_Sorter100|4547_ ;
  assign \new_Sorter100|4647_  = \new_Sorter100|4546_  | \new_Sorter100|4547_ ;
  assign \new_Sorter100|4648_  = \new_Sorter100|4548_  & \new_Sorter100|4549_ ;
  assign \new_Sorter100|4649_  = \new_Sorter100|4548_  | \new_Sorter100|4549_ ;
  assign \new_Sorter100|4650_  = \new_Sorter100|4550_  & \new_Sorter100|4551_ ;
  assign \new_Sorter100|4651_  = \new_Sorter100|4550_  | \new_Sorter100|4551_ ;
  assign \new_Sorter100|4652_  = \new_Sorter100|4552_  & \new_Sorter100|4553_ ;
  assign \new_Sorter100|4653_  = \new_Sorter100|4552_  | \new_Sorter100|4553_ ;
  assign \new_Sorter100|4654_  = \new_Sorter100|4554_  & \new_Sorter100|4555_ ;
  assign \new_Sorter100|4655_  = \new_Sorter100|4554_  | \new_Sorter100|4555_ ;
  assign \new_Sorter100|4656_  = \new_Sorter100|4556_  & \new_Sorter100|4557_ ;
  assign \new_Sorter100|4657_  = \new_Sorter100|4556_  | \new_Sorter100|4557_ ;
  assign \new_Sorter100|4658_  = \new_Sorter100|4558_  & \new_Sorter100|4559_ ;
  assign \new_Sorter100|4659_  = \new_Sorter100|4558_  | \new_Sorter100|4559_ ;
  assign \new_Sorter100|4660_  = \new_Sorter100|4560_  & \new_Sorter100|4561_ ;
  assign \new_Sorter100|4661_  = \new_Sorter100|4560_  | \new_Sorter100|4561_ ;
  assign \new_Sorter100|4662_  = \new_Sorter100|4562_  & \new_Sorter100|4563_ ;
  assign \new_Sorter100|4663_  = \new_Sorter100|4562_  | \new_Sorter100|4563_ ;
  assign \new_Sorter100|4664_  = \new_Sorter100|4564_  & \new_Sorter100|4565_ ;
  assign \new_Sorter100|4665_  = \new_Sorter100|4564_  | \new_Sorter100|4565_ ;
  assign \new_Sorter100|4666_  = \new_Sorter100|4566_  & \new_Sorter100|4567_ ;
  assign \new_Sorter100|4667_  = \new_Sorter100|4566_  | \new_Sorter100|4567_ ;
  assign \new_Sorter100|4668_  = \new_Sorter100|4568_  & \new_Sorter100|4569_ ;
  assign \new_Sorter100|4669_  = \new_Sorter100|4568_  | \new_Sorter100|4569_ ;
  assign \new_Sorter100|4670_  = \new_Sorter100|4570_  & \new_Sorter100|4571_ ;
  assign \new_Sorter100|4671_  = \new_Sorter100|4570_  | \new_Sorter100|4571_ ;
  assign \new_Sorter100|4672_  = \new_Sorter100|4572_  & \new_Sorter100|4573_ ;
  assign \new_Sorter100|4673_  = \new_Sorter100|4572_  | \new_Sorter100|4573_ ;
  assign \new_Sorter100|4674_  = \new_Sorter100|4574_  & \new_Sorter100|4575_ ;
  assign \new_Sorter100|4675_  = \new_Sorter100|4574_  | \new_Sorter100|4575_ ;
  assign \new_Sorter100|4676_  = \new_Sorter100|4576_  & \new_Sorter100|4577_ ;
  assign \new_Sorter100|4677_  = \new_Sorter100|4576_  | \new_Sorter100|4577_ ;
  assign \new_Sorter100|4678_  = \new_Sorter100|4578_  & \new_Sorter100|4579_ ;
  assign \new_Sorter100|4679_  = \new_Sorter100|4578_  | \new_Sorter100|4579_ ;
  assign \new_Sorter100|4680_  = \new_Sorter100|4580_  & \new_Sorter100|4581_ ;
  assign \new_Sorter100|4681_  = \new_Sorter100|4580_  | \new_Sorter100|4581_ ;
  assign \new_Sorter100|4682_  = \new_Sorter100|4582_  & \new_Sorter100|4583_ ;
  assign \new_Sorter100|4683_  = \new_Sorter100|4582_  | \new_Sorter100|4583_ ;
  assign \new_Sorter100|4684_  = \new_Sorter100|4584_  & \new_Sorter100|4585_ ;
  assign \new_Sorter100|4685_  = \new_Sorter100|4584_  | \new_Sorter100|4585_ ;
  assign \new_Sorter100|4686_  = \new_Sorter100|4586_  & \new_Sorter100|4587_ ;
  assign \new_Sorter100|4687_  = \new_Sorter100|4586_  | \new_Sorter100|4587_ ;
  assign \new_Sorter100|4688_  = \new_Sorter100|4588_  & \new_Sorter100|4589_ ;
  assign \new_Sorter100|4689_  = \new_Sorter100|4588_  | \new_Sorter100|4589_ ;
  assign \new_Sorter100|4690_  = \new_Sorter100|4590_  & \new_Sorter100|4591_ ;
  assign \new_Sorter100|4691_  = \new_Sorter100|4590_  | \new_Sorter100|4591_ ;
  assign \new_Sorter100|4692_  = \new_Sorter100|4592_  & \new_Sorter100|4593_ ;
  assign \new_Sorter100|4693_  = \new_Sorter100|4592_  | \new_Sorter100|4593_ ;
  assign \new_Sorter100|4694_  = \new_Sorter100|4594_  & \new_Sorter100|4595_ ;
  assign \new_Sorter100|4695_  = \new_Sorter100|4594_  | \new_Sorter100|4595_ ;
  assign \new_Sorter100|4696_  = \new_Sorter100|4596_  & \new_Sorter100|4597_ ;
  assign \new_Sorter100|4697_  = \new_Sorter100|4596_  | \new_Sorter100|4597_ ;
  assign \new_Sorter100|4698_  = \new_Sorter100|4598_  & \new_Sorter100|4599_ ;
  assign \new_Sorter100|4699_  = \new_Sorter100|4598_  | \new_Sorter100|4599_ ;
  assign \new_Sorter100|4700_  = \new_Sorter100|4600_ ;
  assign \new_Sorter100|4799_  = \new_Sorter100|4699_ ;
  assign \new_Sorter100|4701_  = \new_Sorter100|4601_  & \new_Sorter100|4602_ ;
  assign \new_Sorter100|4702_  = \new_Sorter100|4601_  | \new_Sorter100|4602_ ;
  assign \new_Sorter100|4703_  = \new_Sorter100|4603_  & \new_Sorter100|4604_ ;
  assign \new_Sorter100|4704_  = \new_Sorter100|4603_  | \new_Sorter100|4604_ ;
  assign \new_Sorter100|4705_  = \new_Sorter100|4605_  & \new_Sorter100|4606_ ;
  assign \new_Sorter100|4706_  = \new_Sorter100|4605_  | \new_Sorter100|4606_ ;
  assign \new_Sorter100|4707_  = \new_Sorter100|4607_  & \new_Sorter100|4608_ ;
  assign \new_Sorter100|4708_  = \new_Sorter100|4607_  | \new_Sorter100|4608_ ;
  assign \new_Sorter100|4709_  = \new_Sorter100|4609_  & \new_Sorter100|4610_ ;
  assign \new_Sorter100|4710_  = \new_Sorter100|4609_  | \new_Sorter100|4610_ ;
  assign \new_Sorter100|4711_  = \new_Sorter100|4611_  & \new_Sorter100|4612_ ;
  assign \new_Sorter100|4712_  = \new_Sorter100|4611_  | \new_Sorter100|4612_ ;
  assign \new_Sorter100|4713_  = \new_Sorter100|4613_  & \new_Sorter100|4614_ ;
  assign \new_Sorter100|4714_  = \new_Sorter100|4613_  | \new_Sorter100|4614_ ;
  assign \new_Sorter100|4715_  = \new_Sorter100|4615_  & \new_Sorter100|4616_ ;
  assign \new_Sorter100|4716_  = \new_Sorter100|4615_  | \new_Sorter100|4616_ ;
  assign \new_Sorter100|4717_  = \new_Sorter100|4617_  & \new_Sorter100|4618_ ;
  assign \new_Sorter100|4718_  = \new_Sorter100|4617_  | \new_Sorter100|4618_ ;
  assign \new_Sorter100|4719_  = \new_Sorter100|4619_  & \new_Sorter100|4620_ ;
  assign \new_Sorter100|4720_  = \new_Sorter100|4619_  | \new_Sorter100|4620_ ;
  assign \new_Sorter100|4721_  = \new_Sorter100|4621_  & \new_Sorter100|4622_ ;
  assign \new_Sorter100|4722_  = \new_Sorter100|4621_  | \new_Sorter100|4622_ ;
  assign \new_Sorter100|4723_  = \new_Sorter100|4623_  & \new_Sorter100|4624_ ;
  assign \new_Sorter100|4724_  = \new_Sorter100|4623_  | \new_Sorter100|4624_ ;
  assign \new_Sorter100|4725_  = \new_Sorter100|4625_  & \new_Sorter100|4626_ ;
  assign \new_Sorter100|4726_  = \new_Sorter100|4625_  | \new_Sorter100|4626_ ;
  assign \new_Sorter100|4727_  = \new_Sorter100|4627_  & \new_Sorter100|4628_ ;
  assign \new_Sorter100|4728_  = \new_Sorter100|4627_  | \new_Sorter100|4628_ ;
  assign \new_Sorter100|4729_  = \new_Sorter100|4629_  & \new_Sorter100|4630_ ;
  assign \new_Sorter100|4730_  = \new_Sorter100|4629_  | \new_Sorter100|4630_ ;
  assign \new_Sorter100|4731_  = \new_Sorter100|4631_  & \new_Sorter100|4632_ ;
  assign \new_Sorter100|4732_  = \new_Sorter100|4631_  | \new_Sorter100|4632_ ;
  assign \new_Sorter100|4733_  = \new_Sorter100|4633_  & \new_Sorter100|4634_ ;
  assign \new_Sorter100|4734_  = \new_Sorter100|4633_  | \new_Sorter100|4634_ ;
  assign \new_Sorter100|4735_  = \new_Sorter100|4635_  & \new_Sorter100|4636_ ;
  assign \new_Sorter100|4736_  = \new_Sorter100|4635_  | \new_Sorter100|4636_ ;
  assign \new_Sorter100|4737_  = \new_Sorter100|4637_  & \new_Sorter100|4638_ ;
  assign \new_Sorter100|4738_  = \new_Sorter100|4637_  | \new_Sorter100|4638_ ;
  assign \new_Sorter100|4739_  = \new_Sorter100|4639_  & \new_Sorter100|4640_ ;
  assign \new_Sorter100|4740_  = \new_Sorter100|4639_  | \new_Sorter100|4640_ ;
  assign \new_Sorter100|4741_  = \new_Sorter100|4641_  & \new_Sorter100|4642_ ;
  assign \new_Sorter100|4742_  = \new_Sorter100|4641_  | \new_Sorter100|4642_ ;
  assign \new_Sorter100|4743_  = \new_Sorter100|4643_  & \new_Sorter100|4644_ ;
  assign \new_Sorter100|4744_  = \new_Sorter100|4643_  | \new_Sorter100|4644_ ;
  assign \new_Sorter100|4745_  = \new_Sorter100|4645_  & \new_Sorter100|4646_ ;
  assign \new_Sorter100|4746_  = \new_Sorter100|4645_  | \new_Sorter100|4646_ ;
  assign \new_Sorter100|4747_  = \new_Sorter100|4647_  & \new_Sorter100|4648_ ;
  assign \new_Sorter100|4748_  = \new_Sorter100|4647_  | \new_Sorter100|4648_ ;
  assign \new_Sorter100|4749_  = \new_Sorter100|4649_  & \new_Sorter100|4650_ ;
  assign \new_Sorter100|4750_  = \new_Sorter100|4649_  | \new_Sorter100|4650_ ;
  assign \new_Sorter100|4751_  = \new_Sorter100|4651_  & \new_Sorter100|4652_ ;
  assign \new_Sorter100|4752_  = \new_Sorter100|4651_  | \new_Sorter100|4652_ ;
  assign \new_Sorter100|4753_  = \new_Sorter100|4653_  & \new_Sorter100|4654_ ;
  assign \new_Sorter100|4754_  = \new_Sorter100|4653_  | \new_Sorter100|4654_ ;
  assign \new_Sorter100|4755_  = \new_Sorter100|4655_  & \new_Sorter100|4656_ ;
  assign \new_Sorter100|4756_  = \new_Sorter100|4655_  | \new_Sorter100|4656_ ;
  assign \new_Sorter100|4757_  = \new_Sorter100|4657_  & \new_Sorter100|4658_ ;
  assign \new_Sorter100|4758_  = \new_Sorter100|4657_  | \new_Sorter100|4658_ ;
  assign \new_Sorter100|4759_  = \new_Sorter100|4659_  & \new_Sorter100|4660_ ;
  assign \new_Sorter100|4760_  = \new_Sorter100|4659_  | \new_Sorter100|4660_ ;
  assign \new_Sorter100|4761_  = \new_Sorter100|4661_  & \new_Sorter100|4662_ ;
  assign \new_Sorter100|4762_  = \new_Sorter100|4661_  | \new_Sorter100|4662_ ;
  assign \new_Sorter100|4763_  = \new_Sorter100|4663_  & \new_Sorter100|4664_ ;
  assign \new_Sorter100|4764_  = \new_Sorter100|4663_  | \new_Sorter100|4664_ ;
  assign \new_Sorter100|4765_  = \new_Sorter100|4665_  & \new_Sorter100|4666_ ;
  assign \new_Sorter100|4766_  = \new_Sorter100|4665_  | \new_Sorter100|4666_ ;
  assign \new_Sorter100|4767_  = \new_Sorter100|4667_  & \new_Sorter100|4668_ ;
  assign \new_Sorter100|4768_  = \new_Sorter100|4667_  | \new_Sorter100|4668_ ;
  assign \new_Sorter100|4769_  = \new_Sorter100|4669_  & \new_Sorter100|4670_ ;
  assign \new_Sorter100|4770_  = \new_Sorter100|4669_  | \new_Sorter100|4670_ ;
  assign \new_Sorter100|4771_  = \new_Sorter100|4671_  & \new_Sorter100|4672_ ;
  assign \new_Sorter100|4772_  = \new_Sorter100|4671_  | \new_Sorter100|4672_ ;
  assign \new_Sorter100|4773_  = \new_Sorter100|4673_  & \new_Sorter100|4674_ ;
  assign \new_Sorter100|4774_  = \new_Sorter100|4673_  | \new_Sorter100|4674_ ;
  assign \new_Sorter100|4775_  = \new_Sorter100|4675_  & \new_Sorter100|4676_ ;
  assign \new_Sorter100|4776_  = \new_Sorter100|4675_  | \new_Sorter100|4676_ ;
  assign \new_Sorter100|4777_  = \new_Sorter100|4677_  & \new_Sorter100|4678_ ;
  assign \new_Sorter100|4778_  = \new_Sorter100|4677_  | \new_Sorter100|4678_ ;
  assign \new_Sorter100|4779_  = \new_Sorter100|4679_  & \new_Sorter100|4680_ ;
  assign \new_Sorter100|4780_  = \new_Sorter100|4679_  | \new_Sorter100|4680_ ;
  assign \new_Sorter100|4781_  = \new_Sorter100|4681_  & \new_Sorter100|4682_ ;
  assign \new_Sorter100|4782_  = \new_Sorter100|4681_  | \new_Sorter100|4682_ ;
  assign \new_Sorter100|4783_  = \new_Sorter100|4683_  & \new_Sorter100|4684_ ;
  assign \new_Sorter100|4784_  = \new_Sorter100|4683_  | \new_Sorter100|4684_ ;
  assign \new_Sorter100|4785_  = \new_Sorter100|4685_  & \new_Sorter100|4686_ ;
  assign \new_Sorter100|4786_  = \new_Sorter100|4685_  | \new_Sorter100|4686_ ;
  assign \new_Sorter100|4787_  = \new_Sorter100|4687_  & \new_Sorter100|4688_ ;
  assign \new_Sorter100|4788_  = \new_Sorter100|4687_  | \new_Sorter100|4688_ ;
  assign \new_Sorter100|4789_  = \new_Sorter100|4689_  & \new_Sorter100|4690_ ;
  assign \new_Sorter100|4790_  = \new_Sorter100|4689_  | \new_Sorter100|4690_ ;
  assign \new_Sorter100|4791_  = \new_Sorter100|4691_  & \new_Sorter100|4692_ ;
  assign \new_Sorter100|4792_  = \new_Sorter100|4691_  | \new_Sorter100|4692_ ;
  assign \new_Sorter100|4793_  = \new_Sorter100|4693_  & \new_Sorter100|4694_ ;
  assign \new_Sorter100|4794_  = \new_Sorter100|4693_  | \new_Sorter100|4694_ ;
  assign \new_Sorter100|4795_  = \new_Sorter100|4695_  & \new_Sorter100|4696_ ;
  assign \new_Sorter100|4796_  = \new_Sorter100|4695_  | \new_Sorter100|4696_ ;
  assign \new_Sorter100|4797_  = \new_Sorter100|4697_  & \new_Sorter100|4698_ ;
  assign \new_Sorter100|4798_  = \new_Sorter100|4697_  | \new_Sorter100|4698_ ;
  assign \new_Sorter100|4800_  = \new_Sorter100|4700_  & \new_Sorter100|4701_ ;
  assign \new_Sorter100|4801_  = \new_Sorter100|4700_  | \new_Sorter100|4701_ ;
  assign \new_Sorter100|4802_  = \new_Sorter100|4702_  & \new_Sorter100|4703_ ;
  assign \new_Sorter100|4803_  = \new_Sorter100|4702_  | \new_Sorter100|4703_ ;
  assign \new_Sorter100|4804_  = \new_Sorter100|4704_  & \new_Sorter100|4705_ ;
  assign \new_Sorter100|4805_  = \new_Sorter100|4704_  | \new_Sorter100|4705_ ;
  assign \new_Sorter100|4806_  = \new_Sorter100|4706_  & \new_Sorter100|4707_ ;
  assign \new_Sorter100|4807_  = \new_Sorter100|4706_  | \new_Sorter100|4707_ ;
  assign \new_Sorter100|4808_  = \new_Sorter100|4708_  & \new_Sorter100|4709_ ;
  assign \new_Sorter100|4809_  = \new_Sorter100|4708_  | \new_Sorter100|4709_ ;
  assign \new_Sorter100|4810_  = \new_Sorter100|4710_  & \new_Sorter100|4711_ ;
  assign \new_Sorter100|4811_  = \new_Sorter100|4710_  | \new_Sorter100|4711_ ;
  assign \new_Sorter100|4812_  = \new_Sorter100|4712_  & \new_Sorter100|4713_ ;
  assign \new_Sorter100|4813_  = \new_Sorter100|4712_  | \new_Sorter100|4713_ ;
  assign \new_Sorter100|4814_  = \new_Sorter100|4714_  & \new_Sorter100|4715_ ;
  assign \new_Sorter100|4815_  = \new_Sorter100|4714_  | \new_Sorter100|4715_ ;
  assign \new_Sorter100|4816_  = \new_Sorter100|4716_  & \new_Sorter100|4717_ ;
  assign \new_Sorter100|4817_  = \new_Sorter100|4716_  | \new_Sorter100|4717_ ;
  assign \new_Sorter100|4818_  = \new_Sorter100|4718_  & \new_Sorter100|4719_ ;
  assign \new_Sorter100|4819_  = \new_Sorter100|4718_  | \new_Sorter100|4719_ ;
  assign \new_Sorter100|4820_  = \new_Sorter100|4720_  & \new_Sorter100|4721_ ;
  assign \new_Sorter100|4821_  = \new_Sorter100|4720_  | \new_Sorter100|4721_ ;
  assign \new_Sorter100|4822_  = \new_Sorter100|4722_  & \new_Sorter100|4723_ ;
  assign \new_Sorter100|4823_  = \new_Sorter100|4722_  | \new_Sorter100|4723_ ;
  assign \new_Sorter100|4824_  = \new_Sorter100|4724_  & \new_Sorter100|4725_ ;
  assign \new_Sorter100|4825_  = \new_Sorter100|4724_  | \new_Sorter100|4725_ ;
  assign \new_Sorter100|4826_  = \new_Sorter100|4726_  & \new_Sorter100|4727_ ;
  assign \new_Sorter100|4827_  = \new_Sorter100|4726_  | \new_Sorter100|4727_ ;
  assign \new_Sorter100|4828_  = \new_Sorter100|4728_  & \new_Sorter100|4729_ ;
  assign \new_Sorter100|4829_  = \new_Sorter100|4728_  | \new_Sorter100|4729_ ;
  assign \new_Sorter100|4830_  = \new_Sorter100|4730_  & \new_Sorter100|4731_ ;
  assign \new_Sorter100|4831_  = \new_Sorter100|4730_  | \new_Sorter100|4731_ ;
  assign \new_Sorter100|4832_  = \new_Sorter100|4732_  & \new_Sorter100|4733_ ;
  assign \new_Sorter100|4833_  = \new_Sorter100|4732_  | \new_Sorter100|4733_ ;
  assign \new_Sorter100|4834_  = \new_Sorter100|4734_  & \new_Sorter100|4735_ ;
  assign \new_Sorter100|4835_  = \new_Sorter100|4734_  | \new_Sorter100|4735_ ;
  assign \new_Sorter100|4836_  = \new_Sorter100|4736_  & \new_Sorter100|4737_ ;
  assign \new_Sorter100|4837_  = \new_Sorter100|4736_  | \new_Sorter100|4737_ ;
  assign \new_Sorter100|4838_  = \new_Sorter100|4738_  & \new_Sorter100|4739_ ;
  assign \new_Sorter100|4839_  = \new_Sorter100|4738_  | \new_Sorter100|4739_ ;
  assign \new_Sorter100|4840_  = \new_Sorter100|4740_  & \new_Sorter100|4741_ ;
  assign \new_Sorter100|4841_  = \new_Sorter100|4740_  | \new_Sorter100|4741_ ;
  assign \new_Sorter100|4842_  = \new_Sorter100|4742_  & \new_Sorter100|4743_ ;
  assign \new_Sorter100|4843_  = \new_Sorter100|4742_  | \new_Sorter100|4743_ ;
  assign \new_Sorter100|4844_  = \new_Sorter100|4744_  & \new_Sorter100|4745_ ;
  assign \new_Sorter100|4845_  = \new_Sorter100|4744_  | \new_Sorter100|4745_ ;
  assign \new_Sorter100|4846_  = \new_Sorter100|4746_  & \new_Sorter100|4747_ ;
  assign \new_Sorter100|4847_  = \new_Sorter100|4746_  | \new_Sorter100|4747_ ;
  assign \new_Sorter100|4848_  = \new_Sorter100|4748_  & \new_Sorter100|4749_ ;
  assign \new_Sorter100|4849_  = \new_Sorter100|4748_  | \new_Sorter100|4749_ ;
  assign \new_Sorter100|4850_  = \new_Sorter100|4750_  & \new_Sorter100|4751_ ;
  assign \new_Sorter100|4851_  = \new_Sorter100|4750_  | \new_Sorter100|4751_ ;
  assign \new_Sorter100|4852_  = \new_Sorter100|4752_  & \new_Sorter100|4753_ ;
  assign \new_Sorter100|4853_  = \new_Sorter100|4752_  | \new_Sorter100|4753_ ;
  assign \new_Sorter100|4854_  = \new_Sorter100|4754_  & \new_Sorter100|4755_ ;
  assign \new_Sorter100|4855_  = \new_Sorter100|4754_  | \new_Sorter100|4755_ ;
  assign \new_Sorter100|4856_  = \new_Sorter100|4756_  & \new_Sorter100|4757_ ;
  assign \new_Sorter100|4857_  = \new_Sorter100|4756_  | \new_Sorter100|4757_ ;
  assign \new_Sorter100|4858_  = \new_Sorter100|4758_  & \new_Sorter100|4759_ ;
  assign \new_Sorter100|4859_  = \new_Sorter100|4758_  | \new_Sorter100|4759_ ;
  assign \new_Sorter100|4860_  = \new_Sorter100|4760_  & \new_Sorter100|4761_ ;
  assign \new_Sorter100|4861_  = \new_Sorter100|4760_  | \new_Sorter100|4761_ ;
  assign \new_Sorter100|4862_  = \new_Sorter100|4762_  & \new_Sorter100|4763_ ;
  assign \new_Sorter100|4863_  = \new_Sorter100|4762_  | \new_Sorter100|4763_ ;
  assign \new_Sorter100|4864_  = \new_Sorter100|4764_  & \new_Sorter100|4765_ ;
  assign \new_Sorter100|4865_  = \new_Sorter100|4764_  | \new_Sorter100|4765_ ;
  assign \new_Sorter100|4866_  = \new_Sorter100|4766_  & \new_Sorter100|4767_ ;
  assign \new_Sorter100|4867_  = \new_Sorter100|4766_  | \new_Sorter100|4767_ ;
  assign \new_Sorter100|4868_  = \new_Sorter100|4768_  & \new_Sorter100|4769_ ;
  assign \new_Sorter100|4869_  = \new_Sorter100|4768_  | \new_Sorter100|4769_ ;
  assign \new_Sorter100|4870_  = \new_Sorter100|4770_  & \new_Sorter100|4771_ ;
  assign \new_Sorter100|4871_  = \new_Sorter100|4770_  | \new_Sorter100|4771_ ;
  assign \new_Sorter100|4872_  = \new_Sorter100|4772_  & \new_Sorter100|4773_ ;
  assign \new_Sorter100|4873_  = \new_Sorter100|4772_  | \new_Sorter100|4773_ ;
  assign \new_Sorter100|4874_  = \new_Sorter100|4774_  & \new_Sorter100|4775_ ;
  assign \new_Sorter100|4875_  = \new_Sorter100|4774_  | \new_Sorter100|4775_ ;
  assign \new_Sorter100|4876_  = \new_Sorter100|4776_  & \new_Sorter100|4777_ ;
  assign \new_Sorter100|4877_  = \new_Sorter100|4776_  | \new_Sorter100|4777_ ;
  assign \new_Sorter100|4878_  = \new_Sorter100|4778_  & \new_Sorter100|4779_ ;
  assign \new_Sorter100|4879_  = \new_Sorter100|4778_  | \new_Sorter100|4779_ ;
  assign \new_Sorter100|4880_  = \new_Sorter100|4780_  & \new_Sorter100|4781_ ;
  assign \new_Sorter100|4881_  = \new_Sorter100|4780_  | \new_Sorter100|4781_ ;
  assign \new_Sorter100|4882_  = \new_Sorter100|4782_  & \new_Sorter100|4783_ ;
  assign \new_Sorter100|4883_  = \new_Sorter100|4782_  | \new_Sorter100|4783_ ;
  assign \new_Sorter100|4884_  = \new_Sorter100|4784_  & \new_Sorter100|4785_ ;
  assign \new_Sorter100|4885_  = \new_Sorter100|4784_  | \new_Sorter100|4785_ ;
  assign \new_Sorter100|4886_  = \new_Sorter100|4786_  & \new_Sorter100|4787_ ;
  assign \new_Sorter100|4887_  = \new_Sorter100|4786_  | \new_Sorter100|4787_ ;
  assign \new_Sorter100|4888_  = \new_Sorter100|4788_  & \new_Sorter100|4789_ ;
  assign \new_Sorter100|4889_  = \new_Sorter100|4788_  | \new_Sorter100|4789_ ;
  assign \new_Sorter100|4890_  = \new_Sorter100|4790_  & \new_Sorter100|4791_ ;
  assign \new_Sorter100|4891_  = \new_Sorter100|4790_  | \new_Sorter100|4791_ ;
  assign \new_Sorter100|4892_  = \new_Sorter100|4792_  & \new_Sorter100|4793_ ;
  assign \new_Sorter100|4893_  = \new_Sorter100|4792_  | \new_Sorter100|4793_ ;
  assign \new_Sorter100|4894_  = \new_Sorter100|4794_  & \new_Sorter100|4795_ ;
  assign \new_Sorter100|4895_  = \new_Sorter100|4794_  | \new_Sorter100|4795_ ;
  assign \new_Sorter100|4896_  = \new_Sorter100|4796_  & \new_Sorter100|4797_ ;
  assign \new_Sorter100|4897_  = \new_Sorter100|4796_  | \new_Sorter100|4797_ ;
  assign \new_Sorter100|4898_  = \new_Sorter100|4798_  & \new_Sorter100|4799_ ;
  assign \new_Sorter100|4899_  = \new_Sorter100|4798_  | \new_Sorter100|4799_ ;
  assign \new_Sorter100|4900_  = \new_Sorter100|4800_ ;
  assign \new_Sorter100|4999_  = \new_Sorter100|4899_ ;
  assign \new_Sorter100|4901_  = \new_Sorter100|4801_  & \new_Sorter100|4802_ ;
  assign \new_Sorter100|4902_  = \new_Sorter100|4801_  | \new_Sorter100|4802_ ;
  assign \new_Sorter100|4903_  = \new_Sorter100|4803_  & \new_Sorter100|4804_ ;
  assign \new_Sorter100|4904_  = \new_Sorter100|4803_  | \new_Sorter100|4804_ ;
  assign \new_Sorter100|4905_  = \new_Sorter100|4805_  & \new_Sorter100|4806_ ;
  assign \new_Sorter100|4906_  = \new_Sorter100|4805_  | \new_Sorter100|4806_ ;
  assign \new_Sorter100|4907_  = \new_Sorter100|4807_  & \new_Sorter100|4808_ ;
  assign \new_Sorter100|4908_  = \new_Sorter100|4807_  | \new_Sorter100|4808_ ;
  assign \new_Sorter100|4909_  = \new_Sorter100|4809_  & \new_Sorter100|4810_ ;
  assign \new_Sorter100|4910_  = \new_Sorter100|4809_  | \new_Sorter100|4810_ ;
  assign \new_Sorter100|4911_  = \new_Sorter100|4811_  & \new_Sorter100|4812_ ;
  assign \new_Sorter100|4912_  = \new_Sorter100|4811_  | \new_Sorter100|4812_ ;
  assign \new_Sorter100|4913_  = \new_Sorter100|4813_  & \new_Sorter100|4814_ ;
  assign \new_Sorter100|4914_  = \new_Sorter100|4813_  | \new_Sorter100|4814_ ;
  assign \new_Sorter100|4915_  = \new_Sorter100|4815_  & \new_Sorter100|4816_ ;
  assign \new_Sorter100|4916_  = \new_Sorter100|4815_  | \new_Sorter100|4816_ ;
  assign \new_Sorter100|4917_  = \new_Sorter100|4817_  & \new_Sorter100|4818_ ;
  assign \new_Sorter100|4918_  = \new_Sorter100|4817_  | \new_Sorter100|4818_ ;
  assign \new_Sorter100|4919_  = \new_Sorter100|4819_  & \new_Sorter100|4820_ ;
  assign \new_Sorter100|4920_  = \new_Sorter100|4819_  | \new_Sorter100|4820_ ;
  assign \new_Sorter100|4921_  = \new_Sorter100|4821_  & \new_Sorter100|4822_ ;
  assign \new_Sorter100|4922_  = \new_Sorter100|4821_  | \new_Sorter100|4822_ ;
  assign \new_Sorter100|4923_  = \new_Sorter100|4823_  & \new_Sorter100|4824_ ;
  assign \new_Sorter100|4924_  = \new_Sorter100|4823_  | \new_Sorter100|4824_ ;
  assign \new_Sorter100|4925_  = \new_Sorter100|4825_  & \new_Sorter100|4826_ ;
  assign \new_Sorter100|4926_  = \new_Sorter100|4825_  | \new_Sorter100|4826_ ;
  assign \new_Sorter100|4927_  = \new_Sorter100|4827_  & \new_Sorter100|4828_ ;
  assign \new_Sorter100|4928_  = \new_Sorter100|4827_  | \new_Sorter100|4828_ ;
  assign \new_Sorter100|4929_  = \new_Sorter100|4829_  & \new_Sorter100|4830_ ;
  assign \new_Sorter100|4930_  = \new_Sorter100|4829_  | \new_Sorter100|4830_ ;
  assign \new_Sorter100|4931_  = \new_Sorter100|4831_  & \new_Sorter100|4832_ ;
  assign \new_Sorter100|4932_  = \new_Sorter100|4831_  | \new_Sorter100|4832_ ;
  assign \new_Sorter100|4933_  = \new_Sorter100|4833_  & \new_Sorter100|4834_ ;
  assign \new_Sorter100|4934_  = \new_Sorter100|4833_  | \new_Sorter100|4834_ ;
  assign \new_Sorter100|4935_  = \new_Sorter100|4835_  & \new_Sorter100|4836_ ;
  assign \new_Sorter100|4936_  = \new_Sorter100|4835_  | \new_Sorter100|4836_ ;
  assign \new_Sorter100|4937_  = \new_Sorter100|4837_  & \new_Sorter100|4838_ ;
  assign \new_Sorter100|4938_  = \new_Sorter100|4837_  | \new_Sorter100|4838_ ;
  assign \new_Sorter100|4939_  = \new_Sorter100|4839_  & \new_Sorter100|4840_ ;
  assign \new_Sorter100|4940_  = \new_Sorter100|4839_  | \new_Sorter100|4840_ ;
  assign \new_Sorter100|4941_  = \new_Sorter100|4841_  & \new_Sorter100|4842_ ;
  assign \new_Sorter100|4942_  = \new_Sorter100|4841_  | \new_Sorter100|4842_ ;
  assign \new_Sorter100|4943_  = \new_Sorter100|4843_  & \new_Sorter100|4844_ ;
  assign \new_Sorter100|4944_  = \new_Sorter100|4843_  | \new_Sorter100|4844_ ;
  assign \new_Sorter100|4945_  = \new_Sorter100|4845_  & \new_Sorter100|4846_ ;
  assign \new_Sorter100|4946_  = \new_Sorter100|4845_  | \new_Sorter100|4846_ ;
  assign \new_Sorter100|4947_  = \new_Sorter100|4847_  & \new_Sorter100|4848_ ;
  assign \new_Sorter100|4948_  = \new_Sorter100|4847_  | \new_Sorter100|4848_ ;
  assign \new_Sorter100|4949_  = \new_Sorter100|4849_  & \new_Sorter100|4850_ ;
  assign \new_Sorter100|4950_  = \new_Sorter100|4849_  | \new_Sorter100|4850_ ;
  assign \new_Sorter100|4951_  = \new_Sorter100|4851_  & \new_Sorter100|4852_ ;
  assign \new_Sorter100|4952_  = \new_Sorter100|4851_  | \new_Sorter100|4852_ ;
  assign \new_Sorter100|4953_  = \new_Sorter100|4853_  & \new_Sorter100|4854_ ;
  assign \new_Sorter100|4954_  = \new_Sorter100|4853_  | \new_Sorter100|4854_ ;
  assign \new_Sorter100|4955_  = \new_Sorter100|4855_  & \new_Sorter100|4856_ ;
  assign \new_Sorter100|4956_  = \new_Sorter100|4855_  | \new_Sorter100|4856_ ;
  assign \new_Sorter100|4957_  = \new_Sorter100|4857_  & \new_Sorter100|4858_ ;
  assign \new_Sorter100|4958_  = \new_Sorter100|4857_  | \new_Sorter100|4858_ ;
  assign \new_Sorter100|4959_  = \new_Sorter100|4859_  & \new_Sorter100|4860_ ;
  assign \new_Sorter100|4960_  = \new_Sorter100|4859_  | \new_Sorter100|4860_ ;
  assign \new_Sorter100|4961_  = \new_Sorter100|4861_  & \new_Sorter100|4862_ ;
  assign \new_Sorter100|4962_  = \new_Sorter100|4861_  | \new_Sorter100|4862_ ;
  assign \new_Sorter100|4963_  = \new_Sorter100|4863_  & \new_Sorter100|4864_ ;
  assign \new_Sorter100|4964_  = \new_Sorter100|4863_  | \new_Sorter100|4864_ ;
  assign \new_Sorter100|4965_  = \new_Sorter100|4865_  & \new_Sorter100|4866_ ;
  assign \new_Sorter100|4966_  = \new_Sorter100|4865_  | \new_Sorter100|4866_ ;
  assign \new_Sorter100|4967_  = \new_Sorter100|4867_  & \new_Sorter100|4868_ ;
  assign \new_Sorter100|4968_  = \new_Sorter100|4867_  | \new_Sorter100|4868_ ;
  assign \new_Sorter100|4969_  = \new_Sorter100|4869_  & \new_Sorter100|4870_ ;
  assign \new_Sorter100|4970_  = \new_Sorter100|4869_  | \new_Sorter100|4870_ ;
  assign \new_Sorter100|4971_  = \new_Sorter100|4871_  & \new_Sorter100|4872_ ;
  assign \new_Sorter100|4972_  = \new_Sorter100|4871_  | \new_Sorter100|4872_ ;
  assign \new_Sorter100|4973_  = \new_Sorter100|4873_  & \new_Sorter100|4874_ ;
  assign \new_Sorter100|4974_  = \new_Sorter100|4873_  | \new_Sorter100|4874_ ;
  assign \new_Sorter100|4975_  = \new_Sorter100|4875_  & \new_Sorter100|4876_ ;
  assign \new_Sorter100|4976_  = \new_Sorter100|4875_  | \new_Sorter100|4876_ ;
  assign \new_Sorter100|4977_  = \new_Sorter100|4877_  & \new_Sorter100|4878_ ;
  assign \new_Sorter100|4978_  = \new_Sorter100|4877_  | \new_Sorter100|4878_ ;
  assign \new_Sorter100|4979_  = \new_Sorter100|4879_  & \new_Sorter100|4880_ ;
  assign \new_Sorter100|4980_  = \new_Sorter100|4879_  | \new_Sorter100|4880_ ;
  assign \new_Sorter100|4981_  = \new_Sorter100|4881_  & \new_Sorter100|4882_ ;
  assign \new_Sorter100|4982_  = \new_Sorter100|4881_  | \new_Sorter100|4882_ ;
  assign \new_Sorter100|4983_  = \new_Sorter100|4883_  & \new_Sorter100|4884_ ;
  assign \new_Sorter100|4984_  = \new_Sorter100|4883_  | \new_Sorter100|4884_ ;
  assign \new_Sorter100|4985_  = \new_Sorter100|4885_  & \new_Sorter100|4886_ ;
  assign \new_Sorter100|4986_  = \new_Sorter100|4885_  | \new_Sorter100|4886_ ;
  assign \new_Sorter100|4987_  = \new_Sorter100|4887_  & \new_Sorter100|4888_ ;
  assign \new_Sorter100|4988_  = \new_Sorter100|4887_  | \new_Sorter100|4888_ ;
  assign \new_Sorter100|4989_  = \new_Sorter100|4889_  & \new_Sorter100|4890_ ;
  assign \new_Sorter100|4990_  = \new_Sorter100|4889_  | \new_Sorter100|4890_ ;
  assign \new_Sorter100|4991_  = \new_Sorter100|4891_  & \new_Sorter100|4892_ ;
  assign \new_Sorter100|4992_  = \new_Sorter100|4891_  | \new_Sorter100|4892_ ;
  assign \new_Sorter100|4993_  = \new_Sorter100|4893_  & \new_Sorter100|4894_ ;
  assign \new_Sorter100|4994_  = \new_Sorter100|4893_  | \new_Sorter100|4894_ ;
  assign \new_Sorter100|4995_  = \new_Sorter100|4895_  & \new_Sorter100|4896_ ;
  assign \new_Sorter100|4996_  = \new_Sorter100|4895_  | \new_Sorter100|4896_ ;
  assign \new_Sorter100|4997_  = \new_Sorter100|4897_  & \new_Sorter100|4898_ ;
  assign \new_Sorter100|4998_  = \new_Sorter100|4897_  | \new_Sorter100|4898_ ;
  assign \new_Sorter100|5000_  = \new_Sorter100|4900_  & \new_Sorter100|4901_ ;
  assign \new_Sorter100|5001_  = \new_Sorter100|4900_  | \new_Sorter100|4901_ ;
  assign \new_Sorter100|5002_  = \new_Sorter100|4902_  & \new_Sorter100|4903_ ;
  assign \new_Sorter100|5003_  = \new_Sorter100|4902_  | \new_Sorter100|4903_ ;
  assign \new_Sorter100|5004_  = \new_Sorter100|4904_  & \new_Sorter100|4905_ ;
  assign \new_Sorter100|5005_  = \new_Sorter100|4904_  | \new_Sorter100|4905_ ;
  assign \new_Sorter100|5006_  = \new_Sorter100|4906_  & \new_Sorter100|4907_ ;
  assign \new_Sorter100|5007_  = \new_Sorter100|4906_  | \new_Sorter100|4907_ ;
  assign \new_Sorter100|5008_  = \new_Sorter100|4908_  & \new_Sorter100|4909_ ;
  assign \new_Sorter100|5009_  = \new_Sorter100|4908_  | \new_Sorter100|4909_ ;
  assign \new_Sorter100|5010_  = \new_Sorter100|4910_  & \new_Sorter100|4911_ ;
  assign \new_Sorter100|5011_  = \new_Sorter100|4910_  | \new_Sorter100|4911_ ;
  assign \new_Sorter100|5012_  = \new_Sorter100|4912_  & \new_Sorter100|4913_ ;
  assign \new_Sorter100|5013_  = \new_Sorter100|4912_  | \new_Sorter100|4913_ ;
  assign \new_Sorter100|5014_  = \new_Sorter100|4914_  & \new_Sorter100|4915_ ;
  assign \new_Sorter100|5015_  = \new_Sorter100|4914_  | \new_Sorter100|4915_ ;
  assign \new_Sorter100|5016_  = \new_Sorter100|4916_  & \new_Sorter100|4917_ ;
  assign \new_Sorter100|5017_  = \new_Sorter100|4916_  | \new_Sorter100|4917_ ;
  assign \new_Sorter100|5018_  = \new_Sorter100|4918_  & \new_Sorter100|4919_ ;
  assign \new_Sorter100|5019_  = \new_Sorter100|4918_  | \new_Sorter100|4919_ ;
  assign \new_Sorter100|5020_  = \new_Sorter100|4920_  & \new_Sorter100|4921_ ;
  assign \new_Sorter100|5021_  = \new_Sorter100|4920_  | \new_Sorter100|4921_ ;
  assign \new_Sorter100|5022_  = \new_Sorter100|4922_  & \new_Sorter100|4923_ ;
  assign \new_Sorter100|5023_  = \new_Sorter100|4922_  | \new_Sorter100|4923_ ;
  assign \new_Sorter100|5024_  = \new_Sorter100|4924_  & \new_Sorter100|4925_ ;
  assign \new_Sorter100|5025_  = \new_Sorter100|4924_  | \new_Sorter100|4925_ ;
  assign \new_Sorter100|5026_  = \new_Sorter100|4926_  & \new_Sorter100|4927_ ;
  assign \new_Sorter100|5027_  = \new_Sorter100|4926_  | \new_Sorter100|4927_ ;
  assign \new_Sorter100|5028_  = \new_Sorter100|4928_  & \new_Sorter100|4929_ ;
  assign \new_Sorter100|5029_  = \new_Sorter100|4928_  | \new_Sorter100|4929_ ;
  assign \new_Sorter100|5030_  = \new_Sorter100|4930_  & \new_Sorter100|4931_ ;
  assign \new_Sorter100|5031_  = \new_Sorter100|4930_  | \new_Sorter100|4931_ ;
  assign \new_Sorter100|5032_  = \new_Sorter100|4932_  & \new_Sorter100|4933_ ;
  assign \new_Sorter100|5033_  = \new_Sorter100|4932_  | \new_Sorter100|4933_ ;
  assign \new_Sorter100|5034_  = \new_Sorter100|4934_  & \new_Sorter100|4935_ ;
  assign \new_Sorter100|5035_  = \new_Sorter100|4934_  | \new_Sorter100|4935_ ;
  assign \new_Sorter100|5036_  = \new_Sorter100|4936_  & \new_Sorter100|4937_ ;
  assign \new_Sorter100|5037_  = \new_Sorter100|4936_  | \new_Sorter100|4937_ ;
  assign \new_Sorter100|5038_  = \new_Sorter100|4938_  & \new_Sorter100|4939_ ;
  assign \new_Sorter100|5039_  = \new_Sorter100|4938_  | \new_Sorter100|4939_ ;
  assign \new_Sorter100|5040_  = \new_Sorter100|4940_  & \new_Sorter100|4941_ ;
  assign \new_Sorter100|5041_  = \new_Sorter100|4940_  | \new_Sorter100|4941_ ;
  assign \new_Sorter100|5042_  = \new_Sorter100|4942_  & \new_Sorter100|4943_ ;
  assign \new_Sorter100|5043_  = \new_Sorter100|4942_  | \new_Sorter100|4943_ ;
  assign \new_Sorter100|5044_  = \new_Sorter100|4944_  & \new_Sorter100|4945_ ;
  assign \new_Sorter100|5045_  = \new_Sorter100|4944_  | \new_Sorter100|4945_ ;
  assign \new_Sorter100|5046_  = \new_Sorter100|4946_  & \new_Sorter100|4947_ ;
  assign \new_Sorter100|5047_  = \new_Sorter100|4946_  | \new_Sorter100|4947_ ;
  assign \new_Sorter100|5048_  = \new_Sorter100|4948_  & \new_Sorter100|4949_ ;
  assign \new_Sorter100|5049_  = \new_Sorter100|4948_  | \new_Sorter100|4949_ ;
  assign \new_Sorter100|5050_  = \new_Sorter100|4950_  & \new_Sorter100|4951_ ;
  assign \new_Sorter100|5051_  = \new_Sorter100|4950_  | \new_Sorter100|4951_ ;
  assign \new_Sorter100|5052_  = \new_Sorter100|4952_  & \new_Sorter100|4953_ ;
  assign \new_Sorter100|5053_  = \new_Sorter100|4952_  | \new_Sorter100|4953_ ;
  assign \new_Sorter100|5054_  = \new_Sorter100|4954_  & \new_Sorter100|4955_ ;
  assign \new_Sorter100|5055_  = \new_Sorter100|4954_  | \new_Sorter100|4955_ ;
  assign \new_Sorter100|5056_  = \new_Sorter100|4956_  & \new_Sorter100|4957_ ;
  assign \new_Sorter100|5057_  = \new_Sorter100|4956_  | \new_Sorter100|4957_ ;
  assign \new_Sorter100|5058_  = \new_Sorter100|4958_  & \new_Sorter100|4959_ ;
  assign \new_Sorter100|5059_  = \new_Sorter100|4958_  | \new_Sorter100|4959_ ;
  assign \new_Sorter100|5060_  = \new_Sorter100|4960_  & \new_Sorter100|4961_ ;
  assign \new_Sorter100|5061_  = \new_Sorter100|4960_  | \new_Sorter100|4961_ ;
  assign \new_Sorter100|5062_  = \new_Sorter100|4962_  & \new_Sorter100|4963_ ;
  assign \new_Sorter100|5063_  = \new_Sorter100|4962_  | \new_Sorter100|4963_ ;
  assign \new_Sorter100|5064_  = \new_Sorter100|4964_  & \new_Sorter100|4965_ ;
  assign \new_Sorter100|5065_  = \new_Sorter100|4964_  | \new_Sorter100|4965_ ;
  assign \new_Sorter100|5066_  = \new_Sorter100|4966_  & \new_Sorter100|4967_ ;
  assign \new_Sorter100|5067_  = \new_Sorter100|4966_  | \new_Sorter100|4967_ ;
  assign \new_Sorter100|5068_  = \new_Sorter100|4968_  & \new_Sorter100|4969_ ;
  assign \new_Sorter100|5069_  = \new_Sorter100|4968_  | \new_Sorter100|4969_ ;
  assign \new_Sorter100|5070_  = \new_Sorter100|4970_  & \new_Sorter100|4971_ ;
  assign \new_Sorter100|5071_  = \new_Sorter100|4970_  | \new_Sorter100|4971_ ;
  assign \new_Sorter100|5072_  = \new_Sorter100|4972_  & \new_Sorter100|4973_ ;
  assign \new_Sorter100|5073_  = \new_Sorter100|4972_  | \new_Sorter100|4973_ ;
  assign \new_Sorter100|5074_  = \new_Sorter100|4974_  & \new_Sorter100|4975_ ;
  assign \new_Sorter100|5075_  = \new_Sorter100|4974_  | \new_Sorter100|4975_ ;
  assign \new_Sorter100|5076_  = \new_Sorter100|4976_  & \new_Sorter100|4977_ ;
  assign \new_Sorter100|5077_  = \new_Sorter100|4976_  | \new_Sorter100|4977_ ;
  assign \new_Sorter100|5078_  = \new_Sorter100|4978_  & \new_Sorter100|4979_ ;
  assign \new_Sorter100|5079_  = \new_Sorter100|4978_  | \new_Sorter100|4979_ ;
  assign \new_Sorter100|5080_  = \new_Sorter100|4980_  & \new_Sorter100|4981_ ;
  assign \new_Sorter100|5081_  = \new_Sorter100|4980_  | \new_Sorter100|4981_ ;
  assign \new_Sorter100|5082_  = \new_Sorter100|4982_  & \new_Sorter100|4983_ ;
  assign \new_Sorter100|5083_  = \new_Sorter100|4982_  | \new_Sorter100|4983_ ;
  assign \new_Sorter100|5084_  = \new_Sorter100|4984_  & \new_Sorter100|4985_ ;
  assign \new_Sorter100|5085_  = \new_Sorter100|4984_  | \new_Sorter100|4985_ ;
  assign \new_Sorter100|5086_  = \new_Sorter100|4986_  & \new_Sorter100|4987_ ;
  assign \new_Sorter100|5087_  = \new_Sorter100|4986_  | \new_Sorter100|4987_ ;
  assign \new_Sorter100|5088_  = \new_Sorter100|4988_  & \new_Sorter100|4989_ ;
  assign \new_Sorter100|5089_  = \new_Sorter100|4988_  | \new_Sorter100|4989_ ;
  assign \new_Sorter100|5090_  = \new_Sorter100|4990_  & \new_Sorter100|4991_ ;
  assign \new_Sorter100|5091_  = \new_Sorter100|4990_  | \new_Sorter100|4991_ ;
  assign \new_Sorter100|5092_  = \new_Sorter100|4992_  & \new_Sorter100|4993_ ;
  assign \new_Sorter100|5093_  = \new_Sorter100|4992_  | \new_Sorter100|4993_ ;
  assign \new_Sorter100|5094_  = \new_Sorter100|4994_  & \new_Sorter100|4995_ ;
  assign \new_Sorter100|5095_  = \new_Sorter100|4994_  | \new_Sorter100|4995_ ;
  assign \new_Sorter100|5096_  = \new_Sorter100|4996_  & \new_Sorter100|4997_ ;
  assign \new_Sorter100|5097_  = \new_Sorter100|4996_  | \new_Sorter100|4997_ ;
  assign \new_Sorter100|5098_  = \new_Sorter100|4998_  & \new_Sorter100|4999_ ;
  assign \new_Sorter100|5099_  = \new_Sorter100|4998_  | \new_Sorter100|4999_ ;
  assign \new_Sorter100|5100_  = \new_Sorter100|5000_ ;
  assign \new_Sorter100|5199_  = \new_Sorter100|5099_ ;
  assign \new_Sorter100|5101_  = \new_Sorter100|5001_  & \new_Sorter100|5002_ ;
  assign \new_Sorter100|5102_  = \new_Sorter100|5001_  | \new_Sorter100|5002_ ;
  assign \new_Sorter100|5103_  = \new_Sorter100|5003_  & \new_Sorter100|5004_ ;
  assign \new_Sorter100|5104_  = \new_Sorter100|5003_  | \new_Sorter100|5004_ ;
  assign \new_Sorter100|5105_  = \new_Sorter100|5005_  & \new_Sorter100|5006_ ;
  assign \new_Sorter100|5106_  = \new_Sorter100|5005_  | \new_Sorter100|5006_ ;
  assign \new_Sorter100|5107_  = \new_Sorter100|5007_  & \new_Sorter100|5008_ ;
  assign \new_Sorter100|5108_  = \new_Sorter100|5007_  | \new_Sorter100|5008_ ;
  assign \new_Sorter100|5109_  = \new_Sorter100|5009_  & \new_Sorter100|5010_ ;
  assign \new_Sorter100|5110_  = \new_Sorter100|5009_  | \new_Sorter100|5010_ ;
  assign \new_Sorter100|5111_  = \new_Sorter100|5011_  & \new_Sorter100|5012_ ;
  assign \new_Sorter100|5112_  = \new_Sorter100|5011_  | \new_Sorter100|5012_ ;
  assign \new_Sorter100|5113_  = \new_Sorter100|5013_  & \new_Sorter100|5014_ ;
  assign \new_Sorter100|5114_  = \new_Sorter100|5013_  | \new_Sorter100|5014_ ;
  assign \new_Sorter100|5115_  = \new_Sorter100|5015_  & \new_Sorter100|5016_ ;
  assign \new_Sorter100|5116_  = \new_Sorter100|5015_  | \new_Sorter100|5016_ ;
  assign \new_Sorter100|5117_  = \new_Sorter100|5017_  & \new_Sorter100|5018_ ;
  assign \new_Sorter100|5118_  = \new_Sorter100|5017_  | \new_Sorter100|5018_ ;
  assign \new_Sorter100|5119_  = \new_Sorter100|5019_  & \new_Sorter100|5020_ ;
  assign \new_Sorter100|5120_  = \new_Sorter100|5019_  | \new_Sorter100|5020_ ;
  assign \new_Sorter100|5121_  = \new_Sorter100|5021_  & \new_Sorter100|5022_ ;
  assign \new_Sorter100|5122_  = \new_Sorter100|5021_  | \new_Sorter100|5022_ ;
  assign \new_Sorter100|5123_  = \new_Sorter100|5023_  & \new_Sorter100|5024_ ;
  assign \new_Sorter100|5124_  = \new_Sorter100|5023_  | \new_Sorter100|5024_ ;
  assign \new_Sorter100|5125_  = \new_Sorter100|5025_  & \new_Sorter100|5026_ ;
  assign \new_Sorter100|5126_  = \new_Sorter100|5025_  | \new_Sorter100|5026_ ;
  assign \new_Sorter100|5127_  = \new_Sorter100|5027_  & \new_Sorter100|5028_ ;
  assign \new_Sorter100|5128_  = \new_Sorter100|5027_  | \new_Sorter100|5028_ ;
  assign \new_Sorter100|5129_  = \new_Sorter100|5029_  & \new_Sorter100|5030_ ;
  assign \new_Sorter100|5130_  = \new_Sorter100|5029_  | \new_Sorter100|5030_ ;
  assign \new_Sorter100|5131_  = \new_Sorter100|5031_  & \new_Sorter100|5032_ ;
  assign \new_Sorter100|5132_  = \new_Sorter100|5031_  | \new_Sorter100|5032_ ;
  assign \new_Sorter100|5133_  = \new_Sorter100|5033_  & \new_Sorter100|5034_ ;
  assign \new_Sorter100|5134_  = \new_Sorter100|5033_  | \new_Sorter100|5034_ ;
  assign \new_Sorter100|5135_  = \new_Sorter100|5035_  & \new_Sorter100|5036_ ;
  assign \new_Sorter100|5136_  = \new_Sorter100|5035_  | \new_Sorter100|5036_ ;
  assign \new_Sorter100|5137_  = \new_Sorter100|5037_  & \new_Sorter100|5038_ ;
  assign \new_Sorter100|5138_  = \new_Sorter100|5037_  | \new_Sorter100|5038_ ;
  assign \new_Sorter100|5139_  = \new_Sorter100|5039_  & \new_Sorter100|5040_ ;
  assign \new_Sorter100|5140_  = \new_Sorter100|5039_  | \new_Sorter100|5040_ ;
  assign \new_Sorter100|5141_  = \new_Sorter100|5041_  & \new_Sorter100|5042_ ;
  assign \new_Sorter100|5142_  = \new_Sorter100|5041_  | \new_Sorter100|5042_ ;
  assign \new_Sorter100|5143_  = \new_Sorter100|5043_  & \new_Sorter100|5044_ ;
  assign \new_Sorter100|5144_  = \new_Sorter100|5043_  | \new_Sorter100|5044_ ;
  assign \new_Sorter100|5145_  = \new_Sorter100|5045_  & \new_Sorter100|5046_ ;
  assign \new_Sorter100|5146_  = \new_Sorter100|5045_  | \new_Sorter100|5046_ ;
  assign \new_Sorter100|5147_  = \new_Sorter100|5047_  & \new_Sorter100|5048_ ;
  assign \new_Sorter100|5148_  = \new_Sorter100|5047_  | \new_Sorter100|5048_ ;
  assign \new_Sorter100|5149_  = \new_Sorter100|5049_  & \new_Sorter100|5050_ ;
  assign \new_Sorter100|5150_  = \new_Sorter100|5049_  | \new_Sorter100|5050_ ;
  assign \new_Sorter100|5151_  = \new_Sorter100|5051_  & \new_Sorter100|5052_ ;
  assign \new_Sorter100|5152_  = \new_Sorter100|5051_  | \new_Sorter100|5052_ ;
  assign \new_Sorter100|5153_  = \new_Sorter100|5053_  & \new_Sorter100|5054_ ;
  assign \new_Sorter100|5154_  = \new_Sorter100|5053_  | \new_Sorter100|5054_ ;
  assign \new_Sorter100|5155_  = \new_Sorter100|5055_  & \new_Sorter100|5056_ ;
  assign \new_Sorter100|5156_  = \new_Sorter100|5055_  | \new_Sorter100|5056_ ;
  assign \new_Sorter100|5157_  = \new_Sorter100|5057_  & \new_Sorter100|5058_ ;
  assign \new_Sorter100|5158_  = \new_Sorter100|5057_  | \new_Sorter100|5058_ ;
  assign \new_Sorter100|5159_  = \new_Sorter100|5059_  & \new_Sorter100|5060_ ;
  assign \new_Sorter100|5160_  = \new_Sorter100|5059_  | \new_Sorter100|5060_ ;
  assign \new_Sorter100|5161_  = \new_Sorter100|5061_  & \new_Sorter100|5062_ ;
  assign \new_Sorter100|5162_  = \new_Sorter100|5061_  | \new_Sorter100|5062_ ;
  assign \new_Sorter100|5163_  = \new_Sorter100|5063_  & \new_Sorter100|5064_ ;
  assign \new_Sorter100|5164_  = \new_Sorter100|5063_  | \new_Sorter100|5064_ ;
  assign \new_Sorter100|5165_  = \new_Sorter100|5065_  & \new_Sorter100|5066_ ;
  assign \new_Sorter100|5166_  = \new_Sorter100|5065_  | \new_Sorter100|5066_ ;
  assign \new_Sorter100|5167_  = \new_Sorter100|5067_  & \new_Sorter100|5068_ ;
  assign \new_Sorter100|5168_  = \new_Sorter100|5067_  | \new_Sorter100|5068_ ;
  assign \new_Sorter100|5169_  = \new_Sorter100|5069_  & \new_Sorter100|5070_ ;
  assign \new_Sorter100|5170_  = \new_Sorter100|5069_  | \new_Sorter100|5070_ ;
  assign \new_Sorter100|5171_  = \new_Sorter100|5071_  & \new_Sorter100|5072_ ;
  assign \new_Sorter100|5172_  = \new_Sorter100|5071_  | \new_Sorter100|5072_ ;
  assign \new_Sorter100|5173_  = \new_Sorter100|5073_  & \new_Sorter100|5074_ ;
  assign \new_Sorter100|5174_  = \new_Sorter100|5073_  | \new_Sorter100|5074_ ;
  assign \new_Sorter100|5175_  = \new_Sorter100|5075_  & \new_Sorter100|5076_ ;
  assign \new_Sorter100|5176_  = \new_Sorter100|5075_  | \new_Sorter100|5076_ ;
  assign \new_Sorter100|5177_  = \new_Sorter100|5077_  & \new_Sorter100|5078_ ;
  assign \new_Sorter100|5178_  = \new_Sorter100|5077_  | \new_Sorter100|5078_ ;
  assign \new_Sorter100|5179_  = \new_Sorter100|5079_  & \new_Sorter100|5080_ ;
  assign \new_Sorter100|5180_  = \new_Sorter100|5079_  | \new_Sorter100|5080_ ;
  assign \new_Sorter100|5181_  = \new_Sorter100|5081_  & \new_Sorter100|5082_ ;
  assign \new_Sorter100|5182_  = \new_Sorter100|5081_  | \new_Sorter100|5082_ ;
  assign \new_Sorter100|5183_  = \new_Sorter100|5083_  & \new_Sorter100|5084_ ;
  assign \new_Sorter100|5184_  = \new_Sorter100|5083_  | \new_Sorter100|5084_ ;
  assign \new_Sorter100|5185_  = \new_Sorter100|5085_  & \new_Sorter100|5086_ ;
  assign \new_Sorter100|5186_  = \new_Sorter100|5085_  | \new_Sorter100|5086_ ;
  assign \new_Sorter100|5187_  = \new_Sorter100|5087_  & \new_Sorter100|5088_ ;
  assign \new_Sorter100|5188_  = \new_Sorter100|5087_  | \new_Sorter100|5088_ ;
  assign \new_Sorter100|5189_  = \new_Sorter100|5089_  & \new_Sorter100|5090_ ;
  assign \new_Sorter100|5190_  = \new_Sorter100|5089_  | \new_Sorter100|5090_ ;
  assign \new_Sorter100|5191_  = \new_Sorter100|5091_  & \new_Sorter100|5092_ ;
  assign \new_Sorter100|5192_  = \new_Sorter100|5091_  | \new_Sorter100|5092_ ;
  assign \new_Sorter100|5193_  = \new_Sorter100|5093_  & \new_Sorter100|5094_ ;
  assign \new_Sorter100|5194_  = \new_Sorter100|5093_  | \new_Sorter100|5094_ ;
  assign \new_Sorter100|5195_  = \new_Sorter100|5095_  & \new_Sorter100|5096_ ;
  assign \new_Sorter100|5196_  = \new_Sorter100|5095_  | \new_Sorter100|5096_ ;
  assign \new_Sorter100|5197_  = \new_Sorter100|5097_  & \new_Sorter100|5098_ ;
  assign \new_Sorter100|5198_  = \new_Sorter100|5097_  | \new_Sorter100|5098_ ;
  assign \new_Sorter100|5200_  = \new_Sorter100|5100_  & \new_Sorter100|5101_ ;
  assign \new_Sorter100|5201_  = \new_Sorter100|5100_  | \new_Sorter100|5101_ ;
  assign \new_Sorter100|5202_  = \new_Sorter100|5102_  & \new_Sorter100|5103_ ;
  assign \new_Sorter100|5203_  = \new_Sorter100|5102_  | \new_Sorter100|5103_ ;
  assign \new_Sorter100|5204_  = \new_Sorter100|5104_  & \new_Sorter100|5105_ ;
  assign \new_Sorter100|5205_  = \new_Sorter100|5104_  | \new_Sorter100|5105_ ;
  assign \new_Sorter100|5206_  = \new_Sorter100|5106_  & \new_Sorter100|5107_ ;
  assign \new_Sorter100|5207_  = \new_Sorter100|5106_  | \new_Sorter100|5107_ ;
  assign \new_Sorter100|5208_  = \new_Sorter100|5108_  & \new_Sorter100|5109_ ;
  assign \new_Sorter100|5209_  = \new_Sorter100|5108_  | \new_Sorter100|5109_ ;
  assign \new_Sorter100|5210_  = \new_Sorter100|5110_  & \new_Sorter100|5111_ ;
  assign \new_Sorter100|5211_  = \new_Sorter100|5110_  | \new_Sorter100|5111_ ;
  assign \new_Sorter100|5212_  = \new_Sorter100|5112_  & \new_Sorter100|5113_ ;
  assign \new_Sorter100|5213_  = \new_Sorter100|5112_  | \new_Sorter100|5113_ ;
  assign \new_Sorter100|5214_  = \new_Sorter100|5114_  & \new_Sorter100|5115_ ;
  assign \new_Sorter100|5215_  = \new_Sorter100|5114_  | \new_Sorter100|5115_ ;
  assign \new_Sorter100|5216_  = \new_Sorter100|5116_  & \new_Sorter100|5117_ ;
  assign \new_Sorter100|5217_  = \new_Sorter100|5116_  | \new_Sorter100|5117_ ;
  assign \new_Sorter100|5218_  = \new_Sorter100|5118_  & \new_Sorter100|5119_ ;
  assign \new_Sorter100|5219_  = \new_Sorter100|5118_  | \new_Sorter100|5119_ ;
  assign \new_Sorter100|5220_  = \new_Sorter100|5120_  & \new_Sorter100|5121_ ;
  assign \new_Sorter100|5221_  = \new_Sorter100|5120_  | \new_Sorter100|5121_ ;
  assign \new_Sorter100|5222_  = \new_Sorter100|5122_  & \new_Sorter100|5123_ ;
  assign \new_Sorter100|5223_  = \new_Sorter100|5122_  | \new_Sorter100|5123_ ;
  assign \new_Sorter100|5224_  = \new_Sorter100|5124_  & \new_Sorter100|5125_ ;
  assign \new_Sorter100|5225_  = \new_Sorter100|5124_  | \new_Sorter100|5125_ ;
  assign \new_Sorter100|5226_  = \new_Sorter100|5126_  & \new_Sorter100|5127_ ;
  assign \new_Sorter100|5227_  = \new_Sorter100|5126_  | \new_Sorter100|5127_ ;
  assign \new_Sorter100|5228_  = \new_Sorter100|5128_  & \new_Sorter100|5129_ ;
  assign \new_Sorter100|5229_  = \new_Sorter100|5128_  | \new_Sorter100|5129_ ;
  assign \new_Sorter100|5230_  = \new_Sorter100|5130_  & \new_Sorter100|5131_ ;
  assign \new_Sorter100|5231_  = \new_Sorter100|5130_  | \new_Sorter100|5131_ ;
  assign \new_Sorter100|5232_  = \new_Sorter100|5132_  & \new_Sorter100|5133_ ;
  assign \new_Sorter100|5233_  = \new_Sorter100|5132_  | \new_Sorter100|5133_ ;
  assign \new_Sorter100|5234_  = \new_Sorter100|5134_  & \new_Sorter100|5135_ ;
  assign \new_Sorter100|5235_  = \new_Sorter100|5134_  | \new_Sorter100|5135_ ;
  assign \new_Sorter100|5236_  = \new_Sorter100|5136_  & \new_Sorter100|5137_ ;
  assign \new_Sorter100|5237_  = \new_Sorter100|5136_  | \new_Sorter100|5137_ ;
  assign \new_Sorter100|5238_  = \new_Sorter100|5138_  & \new_Sorter100|5139_ ;
  assign \new_Sorter100|5239_  = \new_Sorter100|5138_  | \new_Sorter100|5139_ ;
  assign \new_Sorter100|5240_  = \new_Sorter100|5140_  & \new_Sorter100|5141_ ;
  assign \new_Sorter100|5241_  = \new_Sorter100|5140_  | \new_Sorter100|5141_ ;
  assign \new_Sorter100|5242_  = \new_Sorter100|5142_  & \new_Sorter100|5143_ ;
  assign \new_Sorter100|5243_  = \new_Sorter100|5142_  | \new_Sorter100|5143_ ;
  assign \new_Sorter100|5244_  = \new_Sorter100|5144_  & \new_Sorter100|5145_ ;
  assign \new_Sorter100|5245_  = \new_Sorter100|5144_  | \new_Sorter100|5145_ ;
  assign \new_Sorter100|5246_  = \new_Sorter100|5146_  & \new_Sorter100|5147_ ;
  assign \new_Sorter100|5247_  = \new_Sorter100|5146_  | \new_Sorter100|5147_ ;
  assign \new_Sorter100|5248_  = \new_Sorter100|5148_  & \new_Sorter100|5149_ ;
  assign \new_Sorter100|5249_  = \new_Sorter100|5148_  | \new_Sorter100|5149_ ;
  assign \new_Sorter100|5250_  = \new_Sorter100|5150_  & \new_Sorter100|5151_ ;
  assign \new_Sorter100|5251_  = \new_Sorter100|5150_  | \new_Sorter100|5151_ ;
  assign \new_Sorter100|5252_  = \new_Sorter100|5152_  & \new_Sorter100|5153_ ;
  assign \new_Sorter100|5253_  = \new_Sorter100|5152_  | \new_Sorter100|5153_ ;
  assign \new_Sorter100|5254_  = \new_Sorter100|5154_  & \new_Sorter100|5155_ ;
  assign \new_Sorter100|5255_  = \new_Sorter100|5154_  | \new_Sorter100|5155_ ;
  assign \new_Sorter100|5256_  = \new_Sorter100|5156_  & \new_Sorter100|5157_ ;
  assign \new_Sorter100|5257_  = \new_Sorter100|5156_  | \new_Sorter100|5157_ ;
  assign \new_Sorter100|5258_  = \new_Sorter100|5158_  & \new_Sorter100|5159_ ;
  assign \new_Sorter100|5259_  = \new_Sorter100|5158_  | \new_Sorter100|5159_ ;
  assign \new_Sorter100|5260_  = \new_Sorter100|5160_  & \new_Sorter100|5161_ ;
  assign \new_Sorter100|5261_  = \new_Sorter100|5160_  | \new_Sorter100|5161_ ;
  assign \new_Sorter100|5262_  = \new_Sorter100|5162_  & \new_Sorter100|5163_ ;
  assign \new_Sorter100|5263_  = \new_Sorter100|5162_  | \new_Sorter100|5163_ ;
  assign \new_Sorter100|5264_  = \new_Sorter100|5164_  & \new_Sorter100|5165_ ;
  assign \new_Sorter100|5265_  = \new_Sorter100|5164_  | \new_Sorter100|5165_ ;
  assign \new_Sorter100|5266_  = \new_Sorter100|5166_  & \new_Sorter100|5167_ ;
  assign \new_Sorter100|5267_  = \new_Sorter100|5166_  | \new_Sorter100|5167_ ;
  assign \new_Sorter100|5268_  = \new_Sorter100|5168_  & \new_Sorter100|5169_ ;
  assign \new_Sorter100|5269_  = \new_Sorter100|5168_  | \new_Sorter100|5169_ ;
  assign \new_Sorter100|5270_  = \new_Sorter100|5170_  & \new_Sorter100|5171_ ;
  assign \new_Sorter100|5271_  = \new_Sorter100|5170_  | \new_Sorter100|5171_ ;
  assign \new_Sorter100|5272_  = \new_Sorter100|5172_  & \new_Sorter100|5173_ ;
  assign \new_Sorter100|5273_  = \new_Sorter100|5172_  | \new_Sorter100|5173_ ;
  assign \new_Sorter100|5274_  = \new_Sorter100|5174_  & \new_Sorter100|5175_ ;
  assign \new_Sorter100|5275_  = \new_Sorter100|5174_  | \new_Sorter100|5175_ ;
  assign \new_Sorter100|5276_  = \new_Sorter100|5176_  & \new_Sorter100|5177_ ;
  assign \new_Sorter100|5277_  = \new_Sorter100|5176_  | \new_Sorter100|5177_ ;
  assign \new_Sorter100|5278_  = \new_Sorter100|5178_  & \new_Sorter100|5179_ ;
  assign \new_Sorter100|5279_  = \new_Sorter100|5178_  | \new_Sorter100|5179_ ;
  assign \new_Sorter100|5280_  = \new_Sorter100|5180_  & \new_Sorter100|5181_ ;
  assign \new_Sorter100|5281_  = \new_Sorter100|5180_  | \new_Sorter100|5181_ ;
  assign \new_Sorter100|5282_  = \new_Sorter100|5182_  & \new_Sorter100|5183_ ;
  assign \new_Sorter100|5283_  = \new_Sorter100|5182_  | \new_Sorter100|5183_ ;
  assign \new_Sorter100|5284_  = \new_Sorter100|5184_  & \new_Sorter100|5185_ ;
  assign \new_Sorter100|5285_  = \new_Sorter100|5184_  | \new_Sorter100|5185_ ;
  assign \new_Sorter100|5286_  = \new_Sorter100|5186_  & \new_Sorter100|5187_ ;
  assign \new_Sorter100|5287_  = \new_Sorter100|5186_  | \new_Sorter100|5187_ ;
  assign \new_Sorter100|5288_  = \new_Sorter100|5188_  & \new_Sorter100|5189_ ;
  assign \new_Sorter100|5289_  = \new_Sorter100|5188_  | \new_Sorter100|5189_ ;
  assign \new_Sorter100|5290_  = \new_Sorter100|5190_  & \new_Sorter100|5191_ ;
  assign \new_Sorter100|5291_  = \new_Sorter100|5190_  | \new_Sorter100|5191_ ;
  assign \new_Sorter100|5292_  = \new_Sorter100|5192_  & \new_Sorter100|5193_ ;
  assign \new_Sorter100|5293_  = \new_Sorter100|5192_  | \new_Sorter100|5193_ ;
  assign \new_Sorter100|5294_  = \new_Sorter100|5194_  & \new_Sorter100|5195_ ;
  assign \new_Sorter100|5295_  = \new_Sorter100|5194_  | \new_Sorter100|5195_ ;
  assign \new_Sorter100|5296_  = \new_Sorter100|5196_  & \new_Sorter100|5197_ ;
  assign \new_Sorter100|5297_  = \new_Sorter100|5196_  | \new_Sorter100|5197_ ;
  assign \new_Sorter100|5298_  = \new_Sorter100|5198_  & \new_Sorter100|5199_ ;
  assign \new_Sorter100|5299_  = \new_Sorter100|5198_  | \new_Sorter100|5199_ ;
  assign \new_Sorter100|5300_  = \new_Sorter100|5200_ ;
  assign \new_Sorter100|5399_  = \new_Sorter100|5299_ ;
  assign \new_Sorter100|5301_  = \new_Sorter100|5201_  & \new_Sorter100|5202_ ;
  assign \new_Sorter100|5302_  = \new_Sorter100|5201_  | \new_Sorter100|5202_ ;
  assign \new_Sorter100|5303_  = \new_Sorter100|5203_  & \new_Sorter100|5204_ ;
  assign \new_Sorter100|5304_  = \new_Sorter100|5203_  | \new_Sorter100|5204_ ;
  assign \new_Sorter100|5305_  = \new_Sorter100|5205_  & \new_Sorter100|5206_ ;
  assign \new_Sorter100|5306_  = \new_Sorter100|5205_  | \new_Sorter100|5206_ ;
  assign \new_Sorter100|5307_  = \new_Sorter100|5207_  & \new_Sorter100|5208_ ;
  assign \new_Sorter100|5308_  = \new_Sorter100|5207_  | \new_Sorter100|5208_ ;
  assign \new_Sorter100|5309_  = \new_Sorter100|5209_  & \new_Sorter100|5210_ ;
  assign \new_Sorter100|5310_  = \new_Sorter100|5209_  | \new_Sorter100|5210_ ;
  assign \new_Sorter100|5311_  = \new_Sorter100|5211_  & \new_Sorter100|5212_ ;
  assign \new_Sorter100|5312_  = \new_Sorter100|5211_  | \new_Sorter100|5212_ ;
  assign \new_Sorter100|5313_  = \new_Sorter100|5213_  & \new_Sorter100|5214_ ;
  assign \new_Sorter100|5314_  = \new_Sorter100|5213_  | \new_Sorter100|5214_ ;
  assign \new_Sorter100|5315_  = \new_Sorter100|5215_  & \new_Sorter100|5216_ ;
  assign \new_Sorter100|5316_  = \new_Sorter100|5215_  | \new_Sorter100|5216_ ;
  assign \new_Sorter100|5317_  = \new_Sorter100|5217_  & \new_Sorter100|5218_ ;
  assign \new_Sorter100|5318_  = \new_Sorter100|5217_  | \new_Sorter100|5218_ ;
  assign \new_Sorter100|5319_  = \new_Sorter100|5219_  & \new_Sorter100|5220_ ;
  assign \new_Sorter100|5320_  = \new_Sorter100|5219_  | \new_Sorter100|5220_ ;
  assign \new_Sorter100|5321_  = \new_Sorter100|5221_  & \new_Sorter100|5222_ ;
  assign \new_Sorter100|5322_  = \new_Sorter100|5221_  | \new_Sorter100|5222_ ;
  assign \new_Sorter100|5323_  = \new_Sorter100|5223_  & \new_Sorter100|5224_ ;
  assign \new_Sorter100|5324_  = \new_Sorter100|5223_  | \new_Sorter100|5224_ ;
  assign \new_Sorter100|5325_  = \new_Sorter100|5225_  & \new_Sorter100|5226_ ;
  assign \new_Sorter100|5326_  = \new_Sorter100|5225_  | \new_Sorter100|5226_ ;
  assign \new_Sorter100|5327_  = \new_Sorter100|5227_  & \new_Sorter100|5228_ ;
  assign \new_Sorter100|5328_  = \new_Sorter100|5227_  | \new_Sorter100|5228_ ;
  assign \new_Sorter100|5329_  = \new_Sorter100|5229_  & \new_Sorter100|5230_ ;
  assign \new_Sorter100|5330_  = \new_Sorter100|5229_  | \new_Sorter100|5230_ ;
  assign \new_Sorter100|5331_  = \new_Sorter100|5231_  & \new_Sorter100|5232_ ;
  assign \new_Sorter100|5332_  = \new_Sorter100|5231_  | \new_Sorter100|5232_ ;
  assign \new_Sorter100|5333_  = \new_Sorter100|5233_  & \new_Sorter100|5234_ ;
  assign \new_Sorter100|5334_  = \new_Sorter100|5233_  | \new_Sorter100|5234_ ;
  assign \new_Sorter100|5335_  = \new_Sorter100|5235_  & \new_Sorter100|5236_ ;
  assign \new_Sorter100|5336_  = \new_Sorter100|5235_  | \new_Sorter100|5236_ ;
  assign \new_Sorter100|5337_  = \new_Sorter100|5237_  & \new_Sorter100|5238_ ;
  assign \new_Sorter100|5338_  = \new_Sorter100|5237_  | \new_Sorter100|5238_ ;
  assign \new_Sorter100|5339_  = \new_Sorter100|5239_  & \new_Sorter100|5240_ ;
  assign \new_Sorter100|5340_  = \new_Sorter100|5239_  | \new_Sorter100|5240_ ;
  assign \new_Sorter100|5341_  = \new_Sorter100|5241_  & \new_Sorter100|5242_ ;
  assign \new_Sorter100|5342_  = \new_Sorter100|5241_  | \new_Sorter100|5242_ ;
  assign \new_Sorter100|5343_  = \new_Sorter100|5243_  & \new_Sorter100|5244_ ;
  assign \new_Sorter100|5344_  = \new_Sorter100|5243_  | \new_Sorter100|5244_ ;
  assign \new_Sorter100|5345_  = \new_Sorter100|5245_  & \new_Sorter100|5246_ ;
  assign \new_Sorter100|5346_  = \new_Sorter100|5245_  | \new_Sorter100|5246_ ;
  assign \new_Sorter100|5347_  = \new_Sorter100|5247_  & \new_Sorter100|5248_ ;
  assign \new_Sorter100|5348_  = \new_Sorter100|5247_  | \new_Sorter100|5248_ ;
  assign \new_Sorter100|5349_  = \new_Sorter100|5249_  & \new_Sorter100|5250_ ;
  assign \new_Sorter100|5350_  = \new_Sorter100|5249_  | \new_Sorter100|5250_ ;
  assign \new_Sorter100|5351_  = \new_Sorter100|5251_  & \new_Sorter100|5252_ ;
  assign \new_Sorter100|5352_  = \new_Sorter100|5251_  | \new_Sorter100|5252_ ;
  assign \new_Sorter100|5353_  = \new_Sorter100|5253_  & \new_Sorter100|5254_ ;
  assign \new_Sorter100|5354_  = \new_Sorter100|5253_  | \new_Sorter100|5254_ ;
  assign \new_Sorter100|5355_  = \new_Sorter100|5255_  & \new_Sorter100|5256_ ;
  assign \new_Sorter100|5356_  = \new_Sorter100|5255_  | \new_Sorter100|5256_ ;
  assign \new_Sorter100|5357_  = \new_Sorter100|5257_  & \new_Sorter100|5258_ ;
  assign \new_Sorter100|5358_  = \new_Sorter100|5257_  | \new_Sorter100|5258_ ;
  assign \new_Sorter100|5359_  = \new_Sorter100|5259_  & \new_Sorter100|5260_ ;
  assign \new_Sorter100|5360_  = \new_Sorter100|5259_  | \new_Sorter100|5260_ ;
  assign \new_Sorter100|5361_  = \new_Sorter100|5261_  & \new_Sorter100|5262_ ;
  assign \new_Sorter100|5362_  = \new_Sorter100|5261_  | \new_Sorter100|5262_ ;
  assign \new_Sorter100|5363_  = \new_Sorter100|5263_  & \new_Sorter100|5264_ ;
  assign \new_Sorter100|5364_  = \new_Sorter100|5263_  | \new_Sorter100|5264_ ;
  assign \new_Sorter100|5365_  = \new_Sorter100|5265_  & \new_Sorter100|5266_ ;
  assign \new_Sorter100|5366_  = \new_Sorter100|5265_  | \new_Sorter100|5266_ ;
  assign \new_Sorter100|5367_  = \new_Sorter100|5267_  & \new_Sorter100|5268_ ;
  assign \new_Sorter100|5368_  = \new_Sorter100|5267_  | \new_Sorter100|5268_ ;
  assign \new_Sorter100|5369_  = \new_Sorter100|5269_  & \new_Sorter100|5270_ ;
  assign \new_Sorter100|5370_  = \new_Sorter100|5269_  | \new_Sorter100|5270_ ;
  assign \new_Sorter100|5371_  = \new_Sorter100|5271_  & \new_Sorter100|5272_ ;
  assign \new_Sorter100|5372_  = \new_Sorter100|5271_  | \new_Sorter100|5272_ ;
  assign \new_Sorter100|5373_  = \new_Sorter100|5273_  & \new_Sorter100|5274_ ;
  assign \new_Sorter100|5374_  = \new_Sorter100|5273_  | \new_Sorter100|5274_ ;
  assign \new_Sorter100|5375_  = \new_Sorter100|5275_  & \new_Sorter100|5276_ ;
  assign \new_Sorter100|5376_  = \new_Sorter100|5275_  | \new_Sorter100|5276_ ;
  assign \new_Sorter100|5377_  = \new_Sorter100|5277_  & \new_Sorter100|5278_ ;
  assign \new_Sorter100|5378_  = \new_Sorter100|5277_  | \new_Sorter100|5278_ ;
  assign \new_Sorter100|5379_  = \new_Sorter100|5279_  & \new_Sorter100|5280_ ;
  assign \new_Sorter100|5380_  = \new_Sorter100|5279_  | \new_Sorter100|5280_ ;
  assign \new_Sorter100|5381_  = \new_Sorter100|5281_  & \new_Sorter100|5282_ ;
  assign \new_Sorter100|5382_  = \new_Sorter100|5281_  | \new_Sorter100|5282_ ;
  assign \new_Sorter100|5383_  = \new_Sorter100|5283_  & \new_Sorter100|5284_ ;
  assign \new_Sorter100|5384_  = \new_Sorter100|5283_  | \new_Sorter100|5284_ ;
  assign \new_Sorter100|5385_  = \new_Sorter100|5285_  & \new_Sorter100|5286_ ;
  assign \new_Sorter100|5386_  = \new_Sorter100|5285_  | \new_Sorter100|5286_ ;
  assign \new_Sorter100|5387_  = \new_Sorter100|5287_  & \new_Sorter100|5288_ ;
  assign \new_Sorter100|5388_  = \new_Sorter100|5287_  | \new_Sorter100|5288_ ;
  assign \new_Sorter100|5389_  = \new_Sorter100|5289_  & \new_Sorter100|5290_ ;
  assign \new_Sorter100|5390_  = \new_Sorter100|5289_  | \new_Sorter100|5290_ ;
  assign \new_Sorter100|5391_  = \new_Sorter100|5291_  & \new_Sorter100|5292_ ;
  assign \new_Sorter100|5392_  = \new_Sorter100|5291_  | \new_Sorter100|5292_ ;
  assign \new_Sorter100|5393_  = \new_Sorter100|5293_  & \new_Sorter100|5294_ ;
  assign \new_Sorter100|5394_  = \new_Sorter100|5293_  | \new_Sorter100|5294_ ;
  assign \new_Sorter100|5395_  = \new_Sorter100|5295_  & \new_Sorter100|5296_ ;
  assign \new_Sorter100|5396_  = \new_Sorter100|5295_  | \new_Sorter100|5296_ ;
  assign \new_Sorter100|5397_  = \new_Sorter100|5297_  & \new_Sorter100|5298_ ;
  assign \new_Sorter100|5398_  = \new_Sorter100|5297_  | \new_Sorter100|5298_ ;
  assign \new_Sorter100|5400_  = \new_Sorter100|5300_  & \new_Sorter100|5301_ ;
  assign \new_Sorter100|5401_  = \new_Sorter100|5300_  | \new_Sorter100|5301_ ;
  assign \new_Sorter100|5402_  = \new_Sorter100|5302_  & \new_Sorter100|5303_ ;
  assign \new_Sorter100|5403_  = \new_Sorter100|5302_  | \new_Sorter100|5303_ ;
  assign \new_Sorter100|5404_  = \new_Sorter100|5304_  & \new_Sorter100|5305_ ;
  assign \new_Sorter100|5405_  = \new_Sorter100|5304_  | \new_Sorter100|5305_ ;
  assign \new_Sorter100|5406_  = \new_Sorter100|5306_  & \new_Sorter100|5307_ ;
  assign \new_Sorter100|5407_  = \new_Sorter100|5306_  | \new_Sorter100|5307_ ;
  assign \new_Sorter100|5408_  = \new_Sorter100|5308_  & \new_Sorter100|5309_ ;
  assign \new_Sorter100|5409_  = \new_Sorter100|5308_  | \new_Sorter100|5309_ ;
  assign \new_Sorter100|5410_  = \new_Sorter100|5310_  & \new_Sorter100|5311_ ;
  assign \new_Sorter100|5411_  = \new_Sorter100|5310_  | \new_Sorter100|5311_ ;
  assign \new_Sorter100|5412_  = \new_Sorter100|5312_  & \new_Sorter100|5313_ ;
  assign \new_Sorter100|5413_  = \new_Sorter100|5312_  | \new_Sorter100|5313_ ;
  assign \new_Sorter100|5414_  = \new_Sorter100|5314_  & \new_Sorter100|5315_ ;
  assign \new_Sorter100|5415_  = \new_Sorter100|5314_  | \new_Sorter100|5315_ ;
  assign \new_Sorter100|5416_  = \new_Sorter100|5316_  & \new_Sorter100|5317_ ;
  assign \new_Sorter100|5417_  = \new_Sorter100|5316_  | \new_Sorter100|5317_ ;
  assign \new_Sorter100|5418_  = \new_Sorter100|5318_  & \new_Sorter100|5319_ ;
  assign \new_Sorter100|5419_  = \new_Sorter100|5318_  | \new_Sorter100|5319_ ;
  assign \new_Sorter100|5420_  = \new_Sorter100|5320_  & \new_Sorter100|5321_ ;
  assign \new_Sorter100|5421_  = \new_Sorter100|5320_  | \new_Sorter100|5321_ ;
  assign \new_Sorter100|5422_  = \new_Sorter100|5322_  & \new_Sorter100|5323_ ;
  assign \new_Sorter100|5423_  = \new_Sorter100|5322_  | \new_Sorter100|5323_ ;
  assign \new_Sorter100|5424_  = \new_Sorter100|5324_  & \new_Sorter100|5325_ ;
  assign \new_Sorter100|5425_  = \new_Sorter100|5324_  | \new_Sorter100|5325_ ;
  assign \new_Sorter100|5426_  = \new_Sorter100|5326_  & \new_Sorter100|5327_ ;
  assign \new_Sorter100|5427_  = \new_Sorter100|5326_  | \new_Sorter100|5327_ ;
  assign \new_Sorter100|5428_  = \new_Sorter100|5328_  & \new_Sorter100|5329_ ;
  assign \new_Sorter100|5429_  = \new_Sorter100|5328_  | \new_Sorter100|5329_ ;
  assign \new_Sorter100|5430_  = \new_Sorter100|5330_  & \new_Sorter100|5331_ ;
  assign \new_Sorter100|5431_  = \new_Sorter100|5330_  | \new_Sorter100|5331_ ;
  assign \new_Sorter100|5432_  = \new_Sorter100|5332_  & \new_Sorter100|5333_ ;
  assign \new_Sorter100|5433_  = \new_Sorter100|5332_  | \new_Sorter100|5333_ ;
  assign \new_Sorter100|5434_  = \new_Sorter100|5334_  & \new_Sorter100|5335_ ;
  assign \new_Sorter100|5435_  = \new_Sorter100|5334_  | \new_Sorter100|5335_ ;
  assign \new_Sorter100|5436_  = \new_Sorter100|5336_  & \new_Sorter100|5337_ ;
  assign \new_Sorter100|5437_  = \new_Sorter100|5336_  | \new_Sorter100|5337_ ;
  assign \new_Sorter100|5438_  = \new_Sorter100|5338_  & \new_Sorter100|5339_ ;
  assign \new_Sorter100|5439_  = \new_Sorter100|5338_  | \new_Sorter100|5339_ ;
  assign \new_Sorter100|5440_  = \new_Sorter100|5340_  & \new_Sorter100|5341_ ;
  assign \new_Sorter100|5441_  = \new_Sorter100|5340_  | \new_Sorter100|5341_ ;
  assign \new_Sorter100|5442_  = \new_Sorter100|5342_  & \new_Sorter100|5343_ ;
  assign \new_Sorter100|5443_  = \new_Sorter100|5342_  | \new_Sorter100|5343_ ;
  assign \new_Sorter100|5444_  = \new_Sorter100|5344_  & \new_Sorter100|5345_ ;
  assign \new_Sorter100|5445_  = \new_Sorter100|5344_  | \new_Sorter100|5345_ ;
  assign \new_Sorter100|5446_  = \new_Sorter100|5346_  & \new_Sorter100|5347_ ;
  assign \new_Sorter100|5447_  = \new_Sorter100|5346_  | \new_Sorter100|5347_ ;
  assign \new_Sorter100|5448_  = \new_Sorter100|5348_  & \new_Sorter100|5349_ ;
  assign \new_Sorter100|5449_  = \new_Sorter100|5348_  | \new_Sorter100|5349_ ;
  assign \new_Sorter100|5450_  = \new_Sorter100|5350_  & \new_Sorter100|5351_ ;
  assign \new_Sorter100|5451_  = \new_Sorter100|5350_  | \new_Sorter100|5351_ ;
  assign \new_Sorter100|5452_  = \new_Sorter100|5352_  & \new_Sorter100|5353_ ;
  assign \new_Sorter100|5453_  = \new_Sorter100|5352_  | \new_Sorter100|5353_ ;
  assign \new_Sorter100|5454_  = \new_Sorter100|5354_  & \new_Sorter100|5355_ ;
  assign \new_Sorter100|5455_  = \new_Sorter100|5354_  | \new_Sorter100|5355_ ;
  assign \new_Sorter100|5456_  = \new_Sorter100|5356_  & \new_Sorter100|5357_ ;
  assign \new_Sorter100|5457_  = \new_Sorter100|5356_  | \new_Sorter100|5357_ ;
  assign \new_Sorter100|5458_  = \new_Sorter100|5358_  & \new_Sorter100|5359_ ;
  assign \new_Sorter100|5459_  = \new_Sorter100|5358_  | \new_Sorter100|5359_ ;
  assign \new_Sorter100|5460_  = \new_Sorter100|5360_  & \new_Sorter100|5361_ ;
  assign \new_Sorter100|5461_  = \new_Sorter100|5360_  | \new_Sorter100|5361_ ;
  assign \new_Sorter100|5462_  = \new_Sorter100|5362_  & \new_Sorter100|5363_ ;
  assign \new_Sorter100|5463_  = \new_Sorter100|5362_  | \new_Sorter100|5363_ ;
  assign \new_Sorter100|5464_  = \new_Sorter100|5364_  & \new_Sorter100|5365_ ;
  assign \new_Sorter100|5465_  = \new_Sorter100|5364_  | \new_Sorter100|5365_ ;
  assign \new_Sorter100|5466_  = \new_Sorter100|5366_  & \new_Sorter100|5367_ ;
  assign \new_Sorter100|5467_  = \new_Sorter100|5366_  | \new_Sorter100|5367_ ;
  assign \new_Sorter100|5468_  = \new_Sorter100|5368_  & \new_Sorter100|5369_ ;
  assign \new_Sorter100|5469_  = \new_Sorter100|5368_  | \new_Sorter100|5369_ ;
  assign \new_Sorter100|5470_  = \new_Sorter100|5370_  & \new_Sorter100|5371_ ;
  assign \new_Sorter100|5471_  = \new_Sorter100|5370_  | \new_Sorter100|5371_ ;
  assign \new_Sorter100|5472_  = \new_Sorter100|5372_  & \new_Sorter100|5373_ ;
  assign \new_Sorter100|5473_  = \new_Sorter100|5372_  | \new_Sorter100|5373_ ;
  assign \new_Sorter100|5474_  = \new_Sorter100|5374_  & \new_Sorter100|5375_ ;
  assign \new_Sorter100|5475_  = \new_Sorter100|5374_  | \new_Sorter100|5375_ ;
  assign \new_Sorter100|5476_  = \new_Sorter100|5376_  & \new_Sorter100|5377_ ;
  assign \new_Sorter100|5477_  = \new_Sorter100|5376_  | \new_Sorter100|5377_ ;
  assign \new_Sorter100|5478_  = \new_Sorter100|5378_  & \new_Sorter100|5379_ ;
  assign \new_Sorter100|5479_  = \new_Sorter100|5378_  | \new_Sorter100|5379_ ;
  assign \new_Sorter100|5480_  = \new_Sorter100|5380_  & \new_Sorter100|5381_ ;
  assign \new_Sorter100|5481_  = \new_Sorter100|5380_  | \new_Sorter100|5381_ ;
  assign \new_Sorter100|5482_  = \new_Sorter100|5382_  & \new_Sorter100|5383_ ;
  assign \new_Sorter100|5483_  = \new_Sorter100|5382_  | \new_Sorter100|5383_ ;
  assign \new_Sorter100|5484_  = \new_Sorter100|5384_  & \new_Sorter100|5385_ ;
  assign \new_Sorter100|5485_  = \new_Sorter100|5384_  | \new_Sorter100|5385_ ;
  assign \new_Sorter100|5486_  = \new_Sorter100|5386_  & \new_Sorter100|5387_ ;
  assign \new_Sorter100|5487_  = \new_Sorter100|5386_  | \new_Sorter100|5387_ ;
  assign \new_Sorter100|5488_  = \new_Sorter100|5388_  & \new_Sorter100|5389_ ;
  assign \new_Sorter100|5489_  = \new_Sorter100|5388_  | \new_Sorter100|5389_ ;
  assign \new_Sorter100|5490_  = \new_Sorter100|5390_  & \new_Sorter100|5391_ ;
  assign \new_Sorter100|5491_  = \new_Sorter100|5390_  | \new_Sorter100|5391_ ;
  assign \new_Sorter100|5492_  = \new_Sorter100|5392_  & \new_Sorter100|5393_ ;
  assign \new_Sorter100|5493_  = \new_Sorter100|5392_  | \new_Sorter100|5393_ ;
  assign \new_Sorter100|5494_  = \new_Sorter100|5394_  & \new_Sorter100|5395_ ;
  assign \new_Sorter100|5495_  = \new_Sorter100|5394_  | \new_Sorter100|5395_ ;
  assign \new_Sorter100|5496_  = \new_Sorter100|5396_  & \new_Sorter100|5397_ ;
  assign \new_Sorter100|5497_  = \new_Sorter100|5396_  | \new_Sorter100|5397_ ;
  assign \new_Sorter100|5498_  = \new_Sorter100|5398_  & \new_Sorter100|5399_ ;
  assign \new_Sorter100|5499_  = \new_Sorter100|5398_  | \new_Sorter100|5399_ ;
  assign \new_Sorter100|5500_  = \new_Sorter100|5400_ ;
  assign \new_Sorter100|5599_  = \new_Sorter100|5499_ ;
  assign \new_Sorter100|5501_  = \new_Sorter100|5401_  & \new_Sorter100|5402_ ;
  assign \new_Sorter100|5502_  = \new_Sorter100|5401_  | \new_Sorter100|5402_ ;
  assign \new_Sorter100|5503_  = \new_Sorter100|5403_  & \new_Sorter100|5404_ ;
  assign \new_Sorter100|5504_  = \new_Sorter100|5403_  | \new_Sorter100|5404_ ;
  assign \new_Sorter100|5505_  = \new_Sorter100|5405_  & \new_Sorter100|5406_ ;
  assign \new_Sorter100|5506_  = \new_Sorter100|5405_  | \new_Sorter100|5406_ ;
  assign \new_Sorter100|5507_  = \new_Sorter100|5407_  & \new_Sorter100|5408_ ;
  assign \new_Sorter100|5508_  = \new_Sorter100|5407_  | \new_Sorter100|5408_ ;
  assign \new_Sorter100|5509_  = \new_Sorter100|5409_  & \new_Sorter100|5410_ ;
  assign \new_Sorter100|5510_  = \new_Sorter100|5409_  | \new_Sorter100|5410_ ;
  assign \new_Sorter100|5511_  = \new_Sorter100|5411_  & \new_Sorter100|5412_ ;
  assign \new_Sorter100|5512_  = \new_Sorter100|5411_  | \new_Sorter100|5412_ ;
  assign \new_Sorter100|5513_  = \new_Sorter100|5413_  & \new_Sorter100|5414_ ;
  assign \new_Sorter100|5514_  = \new_Sorter100|5413_  | \new_Sorter100|5414_ ;
  assign \new_Sorter100|5515_  = \new_Sorter100|5415_  & \new_Sorter100|5416_ ;
  assign \new_Sorter100|5516_  = \new_Sorter100|5415_  | \new_Sorter100|5416_ ;
  assign \new_Sorter100|5517_  = \new_Sorter100|5417_  & \new_Sorter100|5418_ ;
  assign \new_Sorter100|5518_  = \new_Sorter100|5417_  | \new_Sorter100|5418_ ;
  assign \new_Sorter100|5519_  = \new_Sorter100|5419_  & \new_Sorter100|5420_ ;
  assign \new_Sorter100|5520_  = \new_Sorter100|5419_  | \new_Sorter100|5420_ ;
  assign \new_Sorter100|5521_  = \new_Sorter100|5421_  & \new_Sorter100|5422_ ;
  assign \new_Sorter100|5522_  = \new_Sorter100|5421_  | \new_Sorter100|5422_ ;
  assign \new_Sorter100|5523_  = \new_Sorter100|5423_  & \new_Sorter100|5424_ ;
  assign \new_Sorter100|5524_  = \new_Sorter100|5423_  | \new_Sorter100|5424_ ;
  assign \new_Sorter100|5525_  = \new_Sorter100|5425_  & \new_Sorter100|5426_ ;
  assign \new_Sorter100|5526_  = \new_Sorter100|5425_  | \new_Sorter100|5426_ ;
  assign \new_Sorter100|5527_  = \new_Sorter100|5427_  & \new_Sorter100|5428_ ;
  assign \new_Sorter100|5528_  = \new_Sorter100|5427_  | \new_Sorter100|5428_ ;
  assign \new_Sorter100|5529_  = \new_Sorter100|5429_  & \new_Sorter100|5430_ ;
  assign \new_Sorter100|5530_  = \new_Sorter100|5429_  | \new_Sorter100|5430_ ;
  assign \new_Sorter100|5531_  = \new_Sorter100|5431_  & \new_Sorter100|5432_ ;
  assign \new_Sorter100|5532_  = \new_Sorter100|5431_  | \new_Sorter100|5432_ ;
  assign \new_Sorter100|5533_  = \new_Sorter100|5433_  & \new_Sorter100|5434_ ;
  assign \new_Sorter100|5534_  = \new_Sorter100|5433_  | \new_Sorter100|5434_ ;
  assign \new_Sorter100|5535_  = \new_Sorter100|5435_  & \new_Sorter100|5436_ ;
  assign \new_Sorter100|5536_  = \new_Sorter100|5435_  | \new_Sorter100|5436_ ;
  assign \new_Sorter100|5537_  = \new_Sorter100|5437_  & \new_Sorter100|5438_ ;
  assign \new_Sorter100|5538_  = \new_Sorter100|5437_  | \new_Sorter100|5438_ ;
  assign \new_Sorter100|5539_  = \new_Sorter100|5439_  & \new_Sorter100|5440_ ;
  assign \new_Sorter100|5540_  = \new_Sorter100|5439_  | \new_Sorter100|5440_ ;
  assign \new_Sorter100|5541_  = \new_Sorter100|5441_  & \new_Sorter100|5442_ ;
  assign \new_Sorter100|5542_  = \new_Sorter100|5441_  | \new_Sorter100|5442_ ;
  assign \new_Sorter100|5543_  = \new_Sorter100|5443_  & \new_Sorter100|5444_ ;
  assign \new_Sorter100|5544_  = \new_Sorter100|5443_  | \new_Sorter100|5444_ ;
  assign \new_Sorter100|5545_  = \new_Sorter100|5445_  & \new_Sorter100|5446_ ;
  assign \new_Sorter100|5546_  = \new_Sorter100|5445_  | \new_Sorter100|5446_ ;
  assign \new_Sorter100|5547_  = \new_Sorter100|5447_  & \new_Sorter100|5448_ ;
  assign \new_Sorter100|5548_  = \new_Sorter100|5447_  | \new_Sorter100|5448_ ;
  assign \new_Sorter100|5549_  = \new_Sorter100|5449_  & \new_Sorter100|5450_ ;
  assign \new_Sorter100|5550_  = \new_Sorter100|5449_  | \new_Sorter100|5450_ ;
  assign \new_Sorter100|5551_  = \new_Sorter100|5451_  & \new_Sorter100|5452_ ;
  assign \new_Sorter100|5552_  = \new_Sorter100|5451_  | \new_Sorter100|5452_ ;
  assign \new_Sorter100|5553_  = \new_Sorter100|5453_  & \new_Sorter100|5454_ ;
  assign \new_Sorter100|5554_  = \new_Sorter100|5453_  | \new_Sorter100|5454_ ;
  assign \new_Sorter100|5555_  = \new_Sorter100|5455_  & \new_Sorter100|5456_ ;
  assign \new_Sorter100|5556_  = \new_Sorter100|5455_  | \new_Sorter100|5456_ ;
  assign \new_Sorter100|5557_  = \new_Sorter100|5457_  & \new_Sorter100|5458_ ;
  assign \new_Sorter100|5558_  = \new_Sorter100|5457_  | \new_Sorter100|5458_ ;
  assign \new_Sorter100|5559_  = \new_Sorter100|5459_  & \new_Sorter100|5460_ ;
  assign \new_Sorter100|5560_  = \new_Sorter100|5459_  | \new_Sorter100|5460_ ;
  assign \new_Sorter100|5561_  = \new_Sorter100|5461_  & \new_Sorter100|5462_ ;
  assign \new_Sorter100|5562_  = \new_Sorter100|5461_  | \new_Sorter100|5462_ ;
  assign \new_Sorter100|5563_  = \new_Sorter100|5463_  & \new_Sorter100|5464_ ;
  assign \new_Sorter100|5564_  = \new_Sorter100|5463_  | \new_Sorter100|5464_ ;
  assign \new_Sorter100|5565_  = \new_Sorter100|5465_  & \new_Sorter100|5466_ ;
  assign \new_Sorter100|5566_  = \new_Sorter100|5465_  | \new_Sorter100|5466_ ;
  assign \new_Sorter100|5567_  = \new_Sorter100|5467_  & \new_Sorter100|5468_ ;
  assign \new_Sorter100|5568_  = \new_Sorter100|5467_  | \new_Sorter100|5468_ ;
  assign \new_Sorter100|5569_  = \new_Sorter100|5469_  & \new_Sorter100|5470_ ;
  assign \new_Sorter100|5570_  = \new_Sorter100|5469_  | \new_Sorter100|5470_ ;
  assign \new_Sorter100|5571_  = \new_Sorter100|5471_  & \new_Sorter100|5472_ ;
  assign \new_Sorter100|5572_  = \new_Sorter100|5471_  | \new_Sorter100|5472_ ;
  assign \new_Sorter100|5573_  = \new_Sorter100|5473_  & \new_Sorter100|5474_ ;
  assign \new_Sorter100|5574_  = \new_Sorter100|5473_  | \new_Sorter100|5474_ ;
  assign \new_Sorter100|5575_  = \new_Sorter100|5475_  & \new_Sorter100|5476_ ;
  assign \new_Sorter100|5576_  = \new_Sorter100|5475_  | \new_Sorter100|5476_ ;
  assign \new_Sorter100|5577_  = \new_Sorter100|5477_  & \new_Sorter100|5478_ ;
  assign \new_Sorter100|5578_  = \new_Sorter100|5477_  | \new_Sorter100|5478_ ;
  assign \new_Sorter100|5579_  = \new_Sorter100|5479_  & \new_Sorter100|5480_ ;
  assign \new_Sorter100|5580_  = \new_Sorter100|5479_  | \new_Sorter100|5480_ ;
  assign \new_Sorter100|5581_  = \new_Sorter100|5481_  & \new_Sorter100|5482_ ;
  assign \new_Sorter100|5582_  = \new_Sorter100|5481_  | \new_Sorter100|5482_ ;
  assign \new_Sorter100|5583_  = \new_Sorter100|5483_  & \new_Sorter100|5484_ ;
  assign \new_Sorter100|5584_  = \new_Sorter100|5483_  | \new_Sorter100|5484_ ;
  assign \new_Sorter100|5585_  = \new_Sorter100|5485_  & \new_Sorter100|5486_ ;
  assign \new_Sorter100|5586_  = \new_Sorter100|5485_  | \new_Sorter100|5486_ ;
  assign \new_Sorter100|5587_  = \new_Sorter100|5487_  & \new_Sorter100|5488_ ;
  assign \new_Sorter100|5588_  = \new_Sorter100|5487_  | \new_Sorter100|5488_ ;
  assign \new_Sorter100|5589_  = \new_Sorter100|5489_  & \new_Sorter100|5490_ ;
  assign \new_Sorter100|5590_  = \new_Sorter100|5489_  | \new_Sorter100|5490_ ;
  assign \new_Sorter100|5591_  = \new_Sorter100|5491_  & \new_Sorter100|5492_ ;
  assign \new_Sorter100|5592_  = \new_Sorter100|5491_  | \new_Sorter100|5492_ ;
  assign \new_Sorter100|5593_  = \new_Sorter100|5493_  & \new_Sorter100|5494_ ;
  assign \new_Sorter100|5594_  = \new_Sorter100|5493_  | \new_Sorter100|5494_ ;
  assign \new_Sorter100|5595_  = \new_Sorter100|5495_  & \new_Sorter100|5496_ ;
  assign \new_Sorter100|5596_  = \new_Sorter100|5495_  | \new_Sorter100|5496_ ;
  assign \new_Sorter100|5597_  = \new_Sorter100|5497_  & \new_Sorter100|5498_ ;
  assign \new_Sorter100|5598_  = \new_Sorter100|5497_  | \new_Sorter100|5498_ ;
  assign \new_Sorter100|5600_  = \new_Sorter100|5500_  & \new_Sorter100|5501_ ;
  assign \new_Sorter100|5601_  = \new_Sorter100|5500_  | \new_Sorter100|5501_ ;
  assign \new_Sorter100|5602_  = \new_Sorter100|5502_  & \new_Sorter100|5503_ ;
  assign \new_Sorter100|5603_  = \new_Sorter100|5502_  | \new_Sorter100|5503_ ;
  assign \new_Sorter100|5604_  = \new_Sorter100|5504_  & \new_Sorter100|5505_ ;
  assign \new_Sorter100|5605_  = \new_Sorter100|5504_  | \new_Sorter100|5505_ ;
  assign \new_Sorter100|5606_  = \new_Sorter100|5506_  & \new_Sorter100|5507_ ;
  assign \new_Sorter100|5607_  = \new_Sorter100|5506_  | \new_Sorter100|5507_ ;
  assign \new_Sorter100|5608_  = \new_Sorter100|5508_  & \new_Sorter100|5509_ ;
  assign \new_Sorter100|5609_  = \new_Sorter100|5508_  | \new_Sorter100|5509_ ;
  assign \new_Sorter100|5610_  = \new_Sorter100|5510_  & \new_Sorter100|5511_ ;
  assign \new_Sorter100|5611_  = \new_Sorter100|5510_  | \new_Sorter100|5511_ ;
  assign \new_Sorter100|5612_  = \new_Sorter100|5512_  & \new_Sorter100|5513_ ;
  assign \new_Sorter100|5613_  = \new_Sorter100|5512_  | \new_Sorter100|5513_ ;
  assign \new_Sorter100|5614_  = \new_Sorter100|5514_  & \new_Sorter100|5515_ ;
  assign \new_Sorter100|5615_  = \new_Sorter100|5514_  | \new_Sorter100|5515_ ;
  assign \new_Sorter100|5616_  = \new_Sorter100|5516_  & \new_Sorter100|5517_ ;
  assign \new_Sorter100|5617_  = \new_Sorter100|5516_  | \new_Sorter100|5517_ ;
  assign \new_Sorter100|5618_  = \new_Sorter100|5518_  & \new_Sorter100|5519_ ;
  assign \new_Sorter100|5619_  = \new_Sorter100|5518_  | \new_Sorter100|5519_ ;
  assign \new_Sorter100|5620_  = \new_Sorter100|5520_  & \new_Sorter100|5521_ ;
  assign \new_Sorter100|5621_  = \new_Sorter100|5520_  | \new_Sorter100|5521_ ;
  assign \new_Sorter100|5622_  = \new_Sorter100|5522_  & \new_Sorter100|5523_ ;
  assign \new_Sorter100|5623_  = \new_Sorter100|5522_  | \new_Sorter100|5523_ ;
  assign \new_Sorter100|5624_  = \new_Sorter100|5524_  & \new_Sorter100|5525_ ;
  assign \new_Sorter100|5625_  = \new_Sorter100|5524_  | \new_Sorter100|5525_ ;
  assign \new_Sorter100|5626_  = \new_Sorter100|5526_  & \new_Sorter100|5527_ ;
  assign \new_Sorter100|5627_  = \new_Sorter100|5526_  | \new_Sorter100|5527_ ;
  assign \new_Sorter100|5628_  = \new_Sorter100|5528_  & \new_Sorter100|5529_ ;
  assign \new_Sorter100|5629_  = \new_Sorter100|5528_  | \new_Sorter100|5529_ ;
  assign \new_Sorter100|5630_  = \new_Sorter100|5530_  & \new_Sorter100|5531_ ;
  assign \new_Sorter100|5631_  = \new_Sorter100|5530_  | \new_Sorter100|5531_ ;
  assign \new_Sorter100|5632_  = \new_Sorter100|5532_  & \new_Sorter100|5533_ ;
  assign \new_Sorter100|5633_  = \new_Sorter100|5532_  | \new_Sorter100|5533_ ;
  assign \new_Sorter100|5634_  = \new_Sorter100|5534_  & \new_Sorter100|5535_ ;
  assign \new_Sorter100|5635_  = \new_Sorter100|5534_  | \new_Sorter100|5535_ ;
  assign \new_Sorter100|5636_  = \new_Sorter100|5536_  & \new_Sorter100|5537_ ;
  assign \new_Sorter100|5637_  = \new_Sorter100|5536_  | \new_Sorter100|5537_ ;
  assign \new_Sorter100|5638_  = \new_Sorter100|5538_  & \new_Sorter100|5539_ ;
  assign \new_Sorter100|5639_  = \new_Sorter100|5538_  | \new_Sorter100|5539_ ;
  assign \new_Sorter100|5640_  = \new_Sorter100|5540_  & \new_Sorter100|5541_ ;
  assign \new_Sorter100|5641_  = \new_Sorter100|5540_  | \new_Sorter100|5541_ ;
  assign \new_Sorter100|5642_  = \new_Sorter100|5542_  & \new_Sorter100|5543_ ;
  assign \new_Sorter100|5643_  = \new_Sorter100|5542_  | \new_Sorter100|5543_ ;
  assign \new_Sorter100|5644_  = \new_Sorter100|5544_  & \new_Sorter100|5545_ ;
  assign \new_Sorter100|5645_  = \new_Sorter100|5544_  | \new_Sorter100|5545_ ;
  assign \new_Sorter100|5646_  = \new_Sorter100|5546_  & \new_Sorter100|5547_ ;
  assign \new_Sorter100|5647_  = \new_Sorter100|5546_  | \new_Sorter100|5547_ ;
  assign \new_Sorter100|5648_  = \new_Sorter100|5548_  & \new_Sorter100|5549_ ;
  assign \new_Sorter100|5649_  = \new_Sorter100|5548_  | \new_Sorter100|5549_ ;
  assign \new_Sorter100|5650_  = \new_Sorter100|5550_  & \new_Sorter100|5551_ ;
  assign \new_Sorter100|5651_  = \new_Sorter100|5550_  | \new_Sorter100|5551_ ;
  assign \new_Sorter100|5652_  = \new_Sorter100|5552_  & \new_Sorter100|5553_ ;
  assign \new_Sorter100|5653_  = \new_Sorter100|5552_  | \new_Sorter100|5553_ ;
  assign \new_Sorter100|5654_  = \new_Sorter100|5554_  & \new_Sorter100|5555_ ;
  assign \new_Sorter100|5655_  = \new_Sorter100|5554_  | \new_Sorter100|5555_ ;
  assign \new_Sorter100|5656_  = \new_Sorter100|5556_  & \new_Sorter100|5557_ ;
  assign \new_Sorter100|5657_  = \new_Sorter100|5556_  | \new_Sorter100|5557_ ;
  assign \new_Sorter100|5658_  = \new_Sorter100|5558_  & \new_Sorter100|5559_ ;
  assign \new_Sorter100|5659_  = \new_Sorter100|5558_  | \new_Sorter100|5559_ ;
  assign \new_Sorter100|5660_  = \new_Sorter100|5560_  & \new_Sorter100|5561_ ;
  assign \new_Sorter100|5661_  = \new_Sorter100|5560_  | \new_Sorter100|5561_ ;
  assign \new_Sorter100|5662_  = \new_Sorter100|5562_  & \new_Sorter100|5563_ ;
  assign \new_Sorter100|5663_  = \new_Sorter100|5562_  | \new_Sorter100|5563_ ;
  assign \new_Sorter100|5664_  = \new_Sorter100|5564_  & \new_Sorter100|5565_ ;
  assign \new_Sorter100|5665_  = \new_Sorter100|5564_  | \new_Sorter100|5565_ ;
  assign \new_Sorter100|5666_  = \new_Sorter100|5566_  & \new_Sorter100|5567_ ;
  assign \new_Sorter100|5667_  = \new_Sorter100|5566_  | \new_Sorter100|5567_ ;
  assign \new_Sorter100|5668_  = \new_Sorter100|5568_  & \new_Sorter100|5569_ ;
  assign \new_Sorter100|5669_  = \new_Sorter100|5568_  | \new_Sorter100|5569_ ;
  assign \new_Sorter100|5670_  = \new_Sorter100|5570_  & \new_Sorter100|5571_ ;
  assign \new_Sorter100|5671_  = \new_Sorter100|5570_  | \new_Sorter100|5571_ ;
  assign \new_Sorter100|5672_  = \new_Sorter100|5572_  & \new_Sorter100|5573_ ;
  assign \new_Sorter100|5673_  = \new_Sorter100|5572_  | \new_Sorter100|5573_ ;
  assign \new_Sorter100|5674_  = \new_Sorter100|5574_  & \new_Sorter100|5575_ ;
  assign \new_Sorter100|5675_  = \new_Sorter100|5574_  | \new_Sorter100|5575_ ;
  assign \new_Sorter100|5676_  = \new_Sorter100|5576_  & \new_Sorter100|5577_ ;
  assign \new_Sorter100|5677_  = \new_Sorter100|5576_  | \new_Sorter100|5577_ ;
  assign \new_Sorter100|5678_  = \new_Sorter100|5578_  & \new_Sorter100|5579_ ;
  assign \new_Sorter100|5679_  = \new_Sorter100|5578_  | \new_Sorter100|5579_ ;
  assign \new_Sorter100|5680_  = \new_Sorter100|5580_  & \new_Sorter100|5581_ ;
  assign \new_Sorter100|5681_  = \new_Sorter100|5580_  | \new_Sorter100|5581_ ;
  assign \new_Sorter100|5682_  = \new_Sorter100|5582_  & \new_Sorter100|5583_ ;
  assign \new_Sorter100|5683_  = \new_Sorter100|5582_  | \new_Sorter100|5583_ ;
  assign \new_Sorter100|5684_  = \new_Sorter100|5584_  & \new_Sorter100|5585_ ;
  assign \new_Sorter100|5685_  = \new_Sorter100|5584_  | \new_Sorter100|5585_ ;
  assign \new_Sorter100|5686_  = \new_Sorter100|5586_  & \new_Sorter100|5587_ ;
  assign \new_Sorter100|5687_  = \new_Sorter100|5586_  | \new_Sorter100|5587_ ;
  assign \new_Sorter100|5688_  = \new_Sorter100|5588_  & \new_Sorter100|5589_ ;
  assign \new_Sorter100|5689_  = \new_Sorter100|5588_  | \new_Sorter100|5589_ ;
  assign \new_Sorter100|5690_  = \new_Sorter100|5590_  & \new_Sorter100|5591_ ;
  assign \new_Sorter100|5691_  = \new_Sorter100|5590_  | \new_Sorter100|5591_ ;
  assign \new_Sorter100|5692_  = \new_Sorter100|5592_  & \new_Sorter100|5593_ ;
  assign \new_Sorter100|5693_  = \new_Sorter100|5592_  | \new_Sorter100|5593_ ;
  assign \new_Sorter100|5694_  = \new_Sorter100|5594_  & \new_Sorter100|5595_ ;
  assign \new_Sorter100|5695_  = \new_Sorter100|5594_  | \new_Sorter100|5595_ ;
  assign \new_Sorter100|5696_  = \new_Sorter100|5596_  & \new_Sorter100|5597_ ;
  assign \new_Sorter100|5697_  = \new_Sorter100|5596_  | \new_Sorter100|5597_ ;
  assign \new_Sorter100|5698_  = \new_Sorter100|5598_  & \new_Sorter100|5599_ ;
  assign \new_Sorter100|5699_  = \new_Sorter100|5598_  | \new_Sorter100|5599_ ;
  assign \new_Sorter100|5700_  = \new_Sorter100|5600_ ;
  assign \new_Sorter100|5799_  = \new_Sorter100|5699_ ;
  assign \new_Sorter100|5701_  = \new_Sorter100|5601_  & \new_Sorter100|5602_ ;
  assign \new_Sorter100|5702_  = \new_Sorter100|5601_  | \new_Sorter100|5602_ ;
  assign \new_Sorter100|5703_  = \new_Sorter100|5603_  & \new_Sorter100|5604_ ;
  assign \new_Sorter100|5704_  = \new_Sorter100|5603_  | \new_Sorter100|5604_ ;
  assign \new_Sorter100|5705_  = \new_Sorter100|5605_  & \new_Sorter100|5606_ ;
  assign \new_Sorter100|5706_  = \new_Sorter100|5605_  | \new_Sorter100|5606_ ;
  assign \new_Sorter100|5707_  = \new_Sorter100|5607_  & \new_Sorter100|5608_ ;
  assign \new_Sorter100|5708_  = \new_Sorter100|5607_  | \new_Sorter100|5608_ ;
  assign \new_Sorter100|5709_  = \new_Sorter100|5609_  & \new_Sorter100|5610_ ;
  assign \new_Sorter100|5710_  = \new_Sorter100|5609_  | \new_Sorter100|5610_ ;
  assign \new_Sorter100|5711_  = \new_Sorter100|5611_  & \new_Sorter100|5612_ ;
  assign \new_Sorter100|5712_  = \new_Sorter100|5611_  | \new_Sorter100|5612_ ;
  assign \new_Sorter100|5713_  = \new_Sorter100|5613_  & \new_Sorter100|5614_ ;
  assign \new_Sorter100|5714_  = \new_Sorter100|5613_  | \new_Sorter100|5614_ ;
  assign \new_Sorter100|5715_  = \new_Sorter100|5615_  & \new_Sorter100|5616_ ;
  assign \new_Sorter100|5716_  = \new_Sorter100|5615_  | \new_Sorter100|5616_ ;
  assign \new_Sorter100|5717_  = \new_Sorter100|5617_  & \new_Sorter100|5618_ ;
  assign \new_Sorter100|5718_  = \new_Sorter100|5617_  | \new_Sorter100|5618_ ;
  assign \new_Sorter100|5719_  = \new_Sorter100|5619_  & \new_Sorter100|5620_ ;
  assign \new_Sorter100|5720_  = \new_Sorter100|5619_  | \new_Sorter100|5620_ ;
  assign \new_Sorter100|5721_  = \new_Sorter100|5621_  & \new_Sorter100|5622_ ;
  assign \new_Sorter100|5722_  = \new_Sorter100|5621_  | \new_Sorter100|5622_ ;
  assign \new_Sorter100|5723_  = \new_Sorter100|5623_  & \new_Sorter100|5624_ ;
  assign \new_Sorter100|5724_  = \new_Sorter100|5623_  | \new_Sorter100|5624_ ;
  assign \new_Sorter100|5725_  = \new_Sorter100|5625_  & \new_Sorter100|5626_ ;
  assign \new_Sorter100|5726_  = \new_Sorter100|5625_  | \new_Sorter100|5626_ ;
  assign \new_Sorter100|5727_  = \new_Sorter100|5627_  & \new_Sorter100|5628_ ;
  assign \new_Sorter100|5728_  = \new_Sorter100|5627_  | \new_Sorter100|5628_ ;
  assign \new_Sorter100|5729_  = \new_Sorter100|5629_  & \new_Sorter100|5630_ ;
  assign \new_Sorter100|5730_  = \new_Sorter100|5629_  | \new_Sorter100|5630_ ;
  assign \new_Sorter100|5731_  = \new_Sorter100|5631_  & \new_Sorter100|5632_ ;
  assign \new_Sorter100|5732_  = \new_Sorter100|5631_  | \new_Sorter100|5632_ ;
  assign \new_Sorter100|5733_  = \new_Sorter100|5633_  & \new_Sorter100|5634_ ;
  assign \new_Sorter100|5734_  = \new_Sorter100|5633_  | \new_Sorter100|5634_ ;
  assign \new_Sorter100|5735_  = \new_Sorter100|5635_  & \new_Sorter100|5636_ ;
  assign \new_Sorter100|5736_  = \new_Sorter100|5635_  | \new_Sorter100|5636_ ;
  assign \new_Sorter100|5737_  = \new_Sorter100|5637_  & \new_Sorter100|5638_ ;
  assign \new_Sorter100|5738_  = \new_Sorter100|5637_  | \new_Sorter100|5638_ ;
  assign \new_Sorter100|5739_  = \new_Sorter100|5639_  & \new_Sorter100|5640_ ;
  assign \new_Sorter100|5740_  = \new_Sorter100|5639_  | \new_Sorter100|5640_ ;
  assign \new_Sorter100|5741_  = \new_Sorter100|5641_  & \new_Sorter100|5642_ ;
  assign \new_Sorter100|5742_  = \new_Sorter100|5641_  | \new_Sorter100|5642_ ;
  assign \new_Sorter100|5743_  = \new_Sorter100|5643_  & \new_Sorter100|5644_ ;
  assign \new_Sorter100|5744_  = \new_Sorter100|5643_  | \new_Sorter100|5644_ ;
  assign \new_Sorter100|5745_  = \new_Sorter100|5645_  & \new_Sorter100|5646_ ;
  assign \new_Sorter100|5746_  = \new_Sorter100|5645_  | \new_Sorter100|5646_ ;
  assign \new_Sorter100|5747_  = \new_Sorter100|5647_  & \new_Sorter100|5648_ ;
  assign \new_Sorter100|5748_  = \new_Sorter100|5647_  | \new_Sorter100|5648_ ;
  assign \new_Sorter100|5749_  = \new_Sorter100|5649_  & \new_Sorter100|5650_ ;
  assign \new_Sorter100|5750_  = \new_Sorter100|5649_  | \new_Sorter100|5650_ ;
  assign \new_Sorter100|5751_  = \new_Sorter100|5651_  & \new_Sorter100|5652_ ;
  assign \new_Sorter100|5752_  = \new_Sorter100|5651_  | \new_Sorter100|5652_ ;
  assign \new_Sorter100|5753_  = \new_Sorter100|5653_  & \new_Sorter100|5654_ ;
  assign \new_Sorter100|5754_  = \new_Sorter100|5653_  | \new_Sorter100|5654_ ;
  assign \new_Sorter100|5755_  = \new_Sorter100|5655_  & \new_Sorter100|5656_ ;
  assign \new_Sorter100|5756_  = \new_Sorter100|5655_  | \new_Sorter100|5656_ ;
  assign \new_Sorter100|5757_  = \new_Sorter100|5657_  & \new_Sorter100|5658_ ;
  assign \new_Sorter100|5758_  = \new_Sorter100|5657_  | \new_Sorter100|5658_ ;
  assign \new_Sorter100|5759_  = \new_Sorter100|5659_  & \new_Sorter100|5660_ ;
  assign \new_Sorter100|5760_  = \new_Sorter100|5659_  | \new_Sorter100|5660_ ;
  assign \new_Sorter100|5761_  = \new_Sorter100|5661_  & \new_Sorter100|5662_ ;
  assign \new_Sorter100|5762_  = \new_Sorter100|5661_  | \new_Sorter100|5662_ ;
  assign \new_Sorter100|5763_  = \new_Sorter100|5663_  & \new_Sorter100|5664_ ;
  assign \new_Sorter100|5764_  = \new_Sorter100|5663_  | \new_Sorter100|5664_ ;
  assign \new_Sorter100|5765_  = \new_Sorter100|5665_  & \new_Sorter100|5666_ ;
  assign \new_Sorter100|5766_  = \new_Sorter100|5665_  | \new_Sorter100|5666_ ;
  assign \new_Sorter100|5767_  = \new_Sorter100|5667_  & \new_Sorter100|5668_ ;
  assign \new_Sorter100|5768_  = \new_Sorter100|5667_  | \new_Sorter100|5668_ ;
  assign \new_Sorter100|5769_  = \new_Sorter100|5669_  & \new_Sorter100|5670_ ;
  assign \new_Sorter100|5770_  = \new_Sorter100|5669_  | \new_Sorter100|5670_ ;
  assign \new_Sorter100|5771_  = \new_Sorter100|5671_  & \new_Sorter100|5672_ ;
  assign \new_Sorter100|5772_  = \new_Sorter100|5671_  | \new_Sorter100|5672_ ;
  assign \new_Sorter100|5773_  = \new_Sorter100|5673_  & \new_Sorter100|5674_ ;
  assign \new_Sorter100|5774_  = \new_Sorter100|5673_  | \new_Sorter100|5674_ ;
  assign \new_Sorter100|5775_  = \new_Sorter100|5675_  & \new_Sorter100|5676_ ;
  assign \new_Sorter100|5776_  = \new_Sorter100|5675_  | \new_Sorter100|5676_ ;
  assign \new_Sorter100|5777_  = \new_Sorter100|5677_  & \new_Sorter100|5678_ ;
  assign \new_Sorter100|5778_  = \new_Sorter100|5677_  | \new_Sorter100|5678_ ;
  assign \new_Sorter100|5779_  = \new_Sorter100|5679_  & \new_Sorter100|5680_ ;
  assign \new_Sorter100|5780_  = \new_Sorter100|5679_  | \new_Sorter100|5680_ ;
  assign \new_Sorter100|5781_  = \new_Sorter100|5681_  & \new_Sorter100|5682_ ;
  assign \new_Sorter100|5782_  = \new_Sorter100|5681_  | \new_Sorter100|5682_ ;
  assign \new_Sorter100|5783_  = \new_Sorter100|5683_  & \new_Sorter100|5684_ ;
  assign \new_Sorter100|5784_  = \new_Sorter100|5683_  | \new_Sorter100|5684_ ;
  assign \new_Sorter100|5785_  = \new_Sorter100|5685_  & \new_Sorter100|5686_ ;
  assign \new_Sorter100|5786_  = \new_Sorter100|5685_  | \new_Sorter100|5686_ ;
  assign \new_Sorter100|5787_  = \new_Sorter100|5687_  & \new_Sorter100|5688_ ;
  assign \new_Sorter100|5788_  = \new_Sorter100|5687_  | \new_Sorter100|5688_ ;
  assign \new_Sorter100|5789_  = \new_Sorter100|5689_  & \new_Sorter100|5690_ ;
  assign \new_Sorter100|5790_  = \new_Sorter100|5689_  | \new_Sorter100|5690_ ;
  assign \new_Sorter100|5791_  = \new_Sorter100|5691_  & \new_Sorter100|5692_ ;
  assign \new_Sorter100|5792_  = \new_Sorter100|5691_  | \new_Sorter100|5692_ ;
  assign \new_Sorter100|5793_  = \new_Sorter100|5693_  & \new_Sorter100|5694_ ;
  assign \new_Sorter100|5794_  = \new_Sorter100|5693_  | \new_Sorter100|5694_ ;
  assign \new_Sorter100|5795_  = \new_Sorter100|5695_  & \new_Sorter100|5696_ ;
  assign \new_Sorter100|5796_  = \new_Sorter100|5695_  | \new_Sorter100|5696_ ;
  assign \new_Sorter100|5797_  = \new_Sorter100|5697_  & \new_Sorter100|5698_ ;
  assign \new_Sorter100|5798_  = \new_Sorter100|5697_  | \new_Sorter100|5698_ ;
  assign \new_Sorter100|5800_  = \new_Sorter100|5700_  & \new_Sorter100|5701_ ;
  assign \new_Sorter100|5801_  = \new_Sorter100|5700_  | \new_Sorter100|5701_ ;
  assign \new_Sorter100|5802_  = \new_Sorter100|5702_  & \new_Sorter100|5703_ ;
  assign \new_Sorter100|5803_  = \new_Sorter100|5702_  | \new_Sorter100|5703_ ;
  assign \new_Sorter100|5804_  = \new_Sorter100|5704_  & \new_Sorter100|5705_ ;
  assign \new_Sorter100|5805_  = \new_Sorter100|5704_  | \new_Sorter100|5705_ ;
  assign \new_Sorter100|5806_  = \new_Sorter100|5706_  & \new_Sorter100|5707_ ;
  assign \new_Sorter100|5807_  = \new_Sorter100|5706_  | \new_Sorter100|5707_ ;
  assign \new_Sorter100|5808_  = \new_Sorter100|5708_  & \new_Sorter100|5709_ ;
  assign \new_Sorter100|5809_  = \new_Sorter100|5708_  | \new_Sorter100|5709_ ;
  assign \new_Sorter100|5810_  = \new_Sorter100|5710_  & \new_Sorter100|5711_ ;
  assign \new_Sorter100|5811_  = \new_Sorter100|5710_  | \new_Sorter100|5711_ ;
  assign \new_Sorter100|5812_  = \new_Sorter100|5712_  & \new_Sorter100|5713_ ;
  assign \new_Sorter100|5813_  = \new_Sorter100|5712_  | \new_Sorter100|5713_ ;
  assign \new_Sorter100|5814_  = \new_Sorter100|5714_  & \new_Sorter100|5715_ ;
  assign \new_Sorter100|5815_  = \new_Sorter100|5714_  | \new_Sorter100|5715_ ;
  assign \new_Sorter100|5816_  = \new_Sorter100|5716_  & \new_Sorter100|5717_ ;
  assign \new_Sorter100|5817_  = \new_Sorter100|5716_  | \new_Sorter100|5717_ ;
  assign \new_Sorter100|5818_  = \new_Sorter100|5718_  & \new_Sorter100|5719_ ;
  assign \new_Sorter100|5819_  = \new_Sorter100|5718_  | \new_Sorter100|5719_ ;
  assign \new_Sorter100|5820_  = \new_Sorter100|5720_  & \new_Sorter100|5721_ ;
  assign \new_Sorter100|5821_  = \new_Sorter100|5720_  | \new_Sorter100|5721_ ;
  assign \new_Sorter100|5822_  = \new_Sorter100|5722_  & \new_Sorter100|5723_ ;
  assign \new_Sorter100|5823_  = \new_Sorter100|5722_  | \new_Sorter100|5723_ ;
  assign \new_Sorter100|5824_  = \new_Sorter100|5724_  & \new_Sorter100|5725_ ;
  assign \new_Sorter100|5825_  = \new_Sorter100|5724_  | \new_Sorter100|5725_ ;
  assign \new_Sorter100|5826_  = \new_Sorter100|5726_  & \new_Sorter100|5727_ ;
  assign \new_Sorter100|5827_  = \new_Sorter100|5726_  | \new_Sorter100|5727_ ;
  assign \new_Sorter100|5828_  = \new_Sorter100|5728_  & \new_Sorter100|5729_ ;
  assign \new_Sorter100|5829_  = \new_Sorter100|5728_  | \new_Sorter100|5729_ ;
  assign \new_Sorter100|5830_  = \new_Sorter100|5730_  & \new_Sorter100|5731_ ;
  assign \new_Sorter100|5831_  = \new_Sorter100|5730_  | \new_Sorter100|5731_ ;
  assign \new_Sorter100|5832_  = \new_Sorter100|5732_  & \new_Sorter100|5733_ ;
  assign \new_Sorter100|5833_  = \new_Sorter100|5732_  | \new_Sorter100|5733_ ;
  assign \new_Sorter100|5834_  = \new_Sorter100|5734_  & \new_Sorter100|5735_ ;
  assign \new_Sorter100|5835_  = \new_Sorter100|5734_  | \new_Sorter100|5735_ ;
  assign \new_Sorter100|5836_  = \new_Sorter100|5736_  & \new_Sorter100|5737_ ;
  assign \new_Sorter100|5837_  = \new_Sorter100|5736_  | \new_Sorter100|5737_ ;
  assign \new_Sorter100|5838_  = \new_Sorter100|5738_  & \new_Sorter100|5739_ ;
  assign \new_Sorter100|5839_  = \new_Sorter100|5738_  | \new_Sorter100|5739_ ;
  assign \new_Sorter100|5840_  = \new_Sorter100|5740_  & \new_Sorter100|5741_ ;
  assign \new_Sorter100|5841_  = \new_Sorter100|5740_  | \new_Sorter100|5741_ ;
  assign \new_Sorter100|5842_  = \new_Sorter100|5742_  & \new_Sorter100|5743_ ;
  assign \new_Sorter100|5843_  = \new_Sorter100|5742_  | \new_Sorter100|5743_ ;
  assign \new_Sorter100|5844_  = \new_Sorter100|5744_  & \new_Sorter100|5745_ ;
  assign \new_Sorter100|5845_  = \new_Sorter100|5744_  | \new_Sorter100|5745_ ;
  assign \new_Sorter100|5846_  = \new_Sorter100|5746_  & \new_Sorter100|5747_ ;
  assign \new_Sorter100|5847_  = \new_Sorter100|5746_  | \new_Sorter100|5747_ ;
  assign \new_Sorter100|5848_  = \new_Sorter100|5748_  & \new_Sorter100|5749_ ;
  assign \new_Sorter100|5849_  = \new_Sorter100|5748_  | \new_Sorter100|5749_ ;
  assign \new_Sorter100|5850_  = \new_Sorter100|5750_  & \new_Sorter100|5751_ ;
  assign \new_Sorter100|5851_  = \new_Sorter100|5750_  | \new_Sorter100|5751_ ;
  assign \new_Sorter100|5852_  = \new_Sorter100|5752_  & \new_Sorter100|5753_ ;
  assign \new_Sorter100|5853_  = \new_Sorter100|5752_  | \new_Sorter100|5753_ ;
  assign \new_Sorter100|5854_  = \new_Sorter100|5754_  & \new_Sorter100|5755_ ;
  assign \new_Sorter100|5855_  = \new_Sorter100|5754_  | \new_Sorter100|5755_ ;
  assign \new_Sorter100|5856_  = \new_Sorter100|5756_  & \new_Sorter100|5757_ ;
  assign \new_Sorter100|5857_  = \new_Sorter100|5756_  | \new_Sorter100|5757_ ;
  assign \new_Sorter100|5858_  = \new_Sorter100|5758_  & \new_Sorter100|5759_ ;
  assign \new_Sorter100|5859_  = \new_Sorter100|5758_  | \new_Sorter100|5759_ ;
  assign \new_Sorter100|5860_  = \new_Sorter100|5760_  & \new_Sorter100|5761_ ;
  assign \new_Sorter100|5861_  = \new_Sorter100|5760_  | \new_Sorter100|5761_ ;
  assign \new_Sorter100|5862_  = \new_Sorter100|5762_  & \new_Sorter100|5763_ ;
  assign \new_Sorter100|5863_  = \new_Sorter100|5762_  | \new_Sorter100|5763_ ;
  assign \new_Sorter100|5864_  = \new_Sorter100|5764_  & \new_Sorter100|5765_ ;
  assign \new_Sorter100|5865_  = \new_Sorter100|5764_  | \new_Sorter100|5765_ ;
  assign \new_Sorter100|5866_  = \new_Sorter100|5766_  & \new_Sorter100|5767_ ;
  assign \new_Sorter100|5867_  = \new_Sorter100|5766_  | \new_Sorter100|5767_ ;
  assign \new_Sorter100|5868_  = \new_Sorter100|5768_  & \new_Sorter100|5769_ ;
  assign \new_Sorter100|5869_  = \new_Sorter100|5768_  | \new_Sorter100|5769_ ;
  assign \new_Sorter100|5870_  = \new_Sorter100|5770_  & \new_Sorter100|5771_ ;
  assign \new_Sorter100|5871_  = \new_Sorter100|5770_  | \new_Sorter100|5771_ ;
  assign \new_Sorter100|5872_  = \new_Sorter100|5772_  & \new_Sorter100|5773_ ;
  assign \new_Sorter100|5873_  = \new_Sorter100|5772_  | \new_Sorter100|5773_ ;
  assign \new_Sorter100|5874_  = \new_Sorter100|5774_  & \new_Sorter100|5775_ ;
  assign \new_Sorter100|5875_  = \new_Sorter100|5774_  | \new_Sorter100|5775_ ;
  assign \new_Sorter100|5876_  = \new_Sorter100|5776_  & \new_Sorter100|5777_ ;
  assign \new_Sorter100|5877_  = \new_Sorter100|5776_  | \new_Sorter100|5777_ ;
  assign \new_Sorter100|5878_  = \new_Sorter100|5778_  & \new_Sorter100|5779_ ;
  assign \new_Sorter100|5879_  = \new_Sorter100|5778_  | \new_Sorter100|5779_ ;
  assign \new_Sorter100|5880_  = \new_Sorter100|5780_  & \new_Sorter100|5781_ ;
  assign \new_Sorter100|5881_  = \new_Sorter100|5780_  | \new_Sorter100|5781_ ;
  assign \new_Sorter100|5882_  = \new_Sorter100|5782_  & \new_Sorter100|5783_ ;
  assign \new_Sorter100|5883_  = \new_Sorter100|5782_  | \new_Sorter100|5783_ ;
  assign \new_Sorter100|5884_  = \new_Sorter100|5784_  & \new_Sorter100|5785_ ;
  assign \new_Sorter100|5885_  = \new_Sorter100|5784_  | \new_Sorter100|5785_ ;
  assign \new_Sorter100|5886_  = \new_Sorter100|5786_  & \new_Sorter100|5787_ ;
  assign \new_Sorter100|5887_  = \new_Sorter100|5786_  | \new_Sorter100|5787_ ;
  assign \new_Sorter100|5888_  = \new_Sorter100|5788_  & \new_Sorter100|5789_ ;
  assign \new_Sorter100|5889_  = \new_Sorter100|5788_  | \new_Sorter100|5789_ ;
  assign \new_Sorter100|5890_  = \new_Sorter100|5790_  & \new_Sorter100|5791_ ;
  assign \new_Sorter100|5891_  = \new_Sorter100|5790_  | \new_Sorter100|5791_ ;
  assign \new_Sorter100|5892_  = \new_Sorter100|5792_  & \new_Sorter100|5793_ ;
  assign \new_Sorter100|5893_  = \new_Sorter100|5792_  | \new_Sorter100|5793_ ;
  assign \new_Sorter100|5894_  = \new_Sorter100|5794_  & \new_Sorter100|5795_ ;
  assign \new_Sorter100|5895_  = \new_Sorter100|5794_  | \new_Sorter100|5795_ ;
  assign \new_Sorter100|5896_  = \new_Sorter100|5796_  & \new_Sorter100|5797_ ;
  assign \new_Sorter100|5897_  = \new_Sorter100|5796_  | \new_Sorter100|5797_ ;
  assign \new_Sorter100|5898_  = \new_Sorter100|5798_  & \new_Sorter100|5799_ ;
  assign \new_Sorter100|5899_  = \new_Sorter100|5798_  | \new_Sorter100|5799_ ;
  assign \new_Sorter100|5900_  = \new_Sorter100|5800_ ;
  assign \new_Sorter100|5999_  = \new_Sorter100|5899_ ;
  assign \new_Sorter100|5901_  = \new_Sorter100|5801_  & \new_Sorter100|5802_ ;
  assign \new_Sorter100|5902_  = \new_Sorter100|5801_  | \new_Sorter100|5802_ ;
  assign \new_Sorter100|5903_  = \new_Sorter100|5803_  & \new_Sorter100|5804_ ;
  assign \new_Sorter100|5904_  = \new_Sorter100|5803_  | \new_Sorter100|5804_ ;
  assign \new_Sorter100|5905_  = \new_Sorter100|5805_  & \new_Sorter100|5806_ ;
  assign \new_Sorter100|5906_  = \new_Sorter100|5805_  | \new_Sorter100|5806_ ;
  assign \new_Sorter100|5907_  = \new_Sorter100|5807_  & \new_Sorter100|5808_ ;
  assign \new_Sorter100|5908_  = \new_Sorter100|5807_  | \new_Sorter100|5808_ ;
  assign \new_Sorter100|5909_  = \new_Sorter100|5809_  & \new_Sorter100|5810_ ;
  assign \new_Sorter100|5910_  = \new_Sorter100|5809_  | \new_Sorter100|5810_ ;
  assign \new_Sorter100|5911_  = \new_Sorter100|5811_  & \new_Sorter100|5812_ ;
  assign \new_Sorter100|5912_  = \new_Sorter100|5811_  | \new_Sorter100|5812_ ;
  assign \new_Sorter100|5913_  = \new_Sorter100|5813_  & \new_Sorter100|5814_ ;
  assign \new_Sorter100|5914_  = \new_Sorter100|5813_  | \new_Sorter100|5814_ ;
  assign \new_Sorter100|5915_  = \new_Sorter100|5815_  & \new_Sorter100|5816_ ;
  assign \new_Sorter100|5916_  = \new_Sorter100|5815_  | \new_Sorter100|5816_ ;
  assign \new_Sorter100|5917_  = \new_Sorter100|5817_  & \new_Sorter100|5818_ ;
  assign \new_Sorter100|5918_  = \new_Sorter100|5817_  | \new_Sorter100|5818_ ;
  assign \new_Sorter100|5919_  = \new_Sorter100|5819_  & \new_Sorter100|5820_ ;
  assign \new_Sorter100|5920_  = \new_Sorter100|5819_  | \new_Sorter100|5820_ ;
  assign \new_Sorter100|5921_  = \new_Sorter100|5821_  & \new_Sorter100|5822_ ;
  assign \new_Sorter100|5922_  = \new_Sorter100|5821_  | \new_Sorter100|5822_ ;
  assign \new_Sorter100|5923_  = \new_Sorter100|5823_  & \new_Sorter100|5824_ ;
  assign \new_Sorter100|5924_  = \new_Sorter100|5823_  | \new_Sorter100|5824_ ;
  assign \new_Sorter100|5925_  = \new_Sorter100|5825_  & \new_Sorter100|5826_ ;
  assign \new_Sorter100|5926_  = \new_Sorter100|5825_  | \new_Sorter100|5826_ ;
  assign \new_Sorter100|5927_  = \new_Sorter100|5827_  & \new_Sorter100|5828_ ;
  assign \new_Sorter100|5928_  = \new_Sorter100|5827_  | \new_Sorter100|5828_ ;
  assign \new_Sorter100|5929_  = \new_Sorter100|5829_  & \new_Sorter100|5830_ ;
  assign \new_Sorter100|5930_  = \new_Sorter100|5829_  | \new_Sorter100|5830_ ;
  assign \new_Sorter100|5931_  = \new_Sorter100|5831_  & \new_Sorter100|5832_ ;
  assign \new_Sorter100|5932_  = \new_Sorter100|5831_  | \new_Sorter100|5832_ ;
  assign \new_Sorter100|5933_  = \new_Sorter100|5833_  & \new_Sorter100|5834_ ;
  assign \new_Sorter100|5934_  = \new_Sorter100|5833_  | \new_Sorter100|5834_ ;
  assign \new_Sorter100|5935_  = \new_Sorter100|5835_  & \new_Sorter100|5836_ ;
  assign \new_Sorter100|5936_  = \new_Sorter100|5835_  | \new_Sorter100|5836_ ;
  assign \new_Sorter100|5937_  = \new_Sorter100|5837_  & \new_Sorter100|5838_ ;
  assign \new_Sorter100|5938_  = \new_Sorter100|5837_  | \new_Sorter100|5838_ ;
  assign \new_Sorter100|5939_  = \new_Sorter100|5839_  & \new_Sorter100|5840_ ;
  assign \new_Sorter100|5940_  = \new_Sorter100|5839_  | \new_Sorter100|5840_ ;
  assign \new_Sorter100|5941_  = \new_Sorter100|5841_  & \new_Sorter100|5842_ ;
  assign \new_Sorter100|5942_  = \new_Sorter100|5841_  | \new_Sorter100|5842_ ;
  assign \new_Sorter100|5943_  = \new_Sorter100|5843_  & \new_Sorter100|5844_ ;
  assign \new_Sorter100|5944_  = \new_Sorter100|5843_  | \new_Sorter100|5844_ ;
  assign \new_Sorter100|5945_  = \new_Sorter100|5845_  & \new_Sorter100|5846_ ;
  assign \new_Sorter100|5946_  = \new_Sorter100|5845_  | \new_Sorter100|5846_ ;
  assign \new_Sorter100|5947_  = \new_Sorter100|5847_  & \new_Sorter100|5848_ ;
  assign \new_Sorter100|5948_  = \new_Sorter100|5847_  | \new_Sorter100|5848_ ;
  assign \new_Sorter100|5949_  = \new_Sorter100|5849_  & \new_Sorter100|5850_ ;
  assign \new_Sorter100|5950_  = \new_Sorter100|5849_  | \new_Sorter100|5850_ ;
  assign \new_Sorter100|5951_  = \new_Sorter100|5851_  & \new_Sorter100|5852_ ;
  assign \new_Sorter100|5952_  = \new_Sorter100|5851_  | \new_Sorter100|5852_ ;
  assign \new_Sorter100|5953_  = \new_Sorter100|5853_  & \new_Sorter100|5854_ ;
  assign \new_Sorter100|5954_  = \new_Sorter100|5853_  | \new_Sorter100|5854_ ;
  assign \new_Sorter100|5955_  = \new_Sorter100|5855_  & \new_Sorter100|5856_ ;
  assign \new_Sorter100|5956_  = \new_Sorter100|5855_  | \new_Sorter100|5856_ ;
  assign \new_Sorter100|5957_  = \new_Sorter100|5857_  & \new_Sorter100|5858_ ;
  assign \new_Sorter100|5958_  = \new_Sorter100|5857_  | \new_Sorter100|5858_ ;
  assign \new_Sorter100|5959_  = \new_Sorter100|5859_  & \new_Sorter100|5860_ ;
  assign \new_Sorter100|5960_  = \new_Sorter100|5859_  | \new_Sorter100|5860_ ;
  assign \new_Sorter100|5961_  = \new_Sorter100|5861_  & \new_Sorter100|5862_ ;
  assign \new_Sorter100|5962_  = \new_Sorter100|5861_  | \new_Sorter100|5862_ ;
  assign \new_Sorter100|5963_  = \new_Sorter100|5863_  & \new_Sorter100|5864_ ;
  assign \new_Sorter100|5964_  = \new_Sorter100|5863_  | \new_Sorter100|5864_ ;
  assign \new_Sorter100|5965_  = \new_Sorter100|5865_  & \new_Sorter100|5866_ ;
  assign \new_Sorter100|5966_  = \new_Sorter100|5865_  | \new_Sorter100|5866_ ;
  assign \new_Sorter100|5967_  = \new_Sorter100|5867_  & \new_Sorter100|5868_ ;
  assign \new_Sorter100|5968_  = \new_Sorter100|5867_  | \new_Sorter100|5868_ ;
  assign \new_Sorter100|5969_  = \new_Sorter100|5869_  & \new_Sorter100|5870_ ;
  assign \new_Sorter100|5970_  = \new_Sorter100|5869_  | \new_Sorter100|5870_ ;
  assign \new_Sorter100|5971_  = \new_Sorter100|5871_  & \new_Sorter100|5872_ ;
  assign \new_Sorter100|5972_  = \new_Sorter100|5871_  | \new_Sorter100|5872_ ;
  assign \new_Sorter100|5973_  = \new_Sorter100|5873_  & \new_Sorter100|5874_ ;
  assign \new_Sorter100|5974_  = \new_Sorter100|5873_  | \new_Sorter100|5874_ ;
  assign \new_Sorter100|5975_  = \new_Sorter100|5875_  & \new_Sorter100|5876_ ;
  assign \new_Sorter100|5976_  = \new_Sorter100|5875_  | \new_Sorter100|5876_ ;
  assign \new_Sorter100|5977_  = \new_Sorter100|5877_  & \new_Sorter100|5878_ ;
  assign \new_Sorter100|5978_  = \new_Sorter100|5877_  | \new_Sorter100|5878_ ;
  assign \new_Sorter100|5979_  = \new_Sorter100|5879_  & \new_Sorter100|5880_ ;
  assign \new_Sorter100|5980_  = \new_Sorter100|5879_  | \new_Sorter100|5880_ ;
  assign \new_Sorter100|5981_  = \new_Sorter100|5881_  & \new_Sorter100|5882_ ;
  assign \new_Sorter100|5982_  = \new_Sorter100|5881_  | \new_Sorter100|5882_ ;
  assign \new_Sorter100|5983_  = \new_Sorter100|5883_  & \new_Sorter100|5884_ ;
  assign \new_Sorter100|5984_  = \new_Sorter100|5883_  | \new_Sorter100|5884_ ;
  assign \new_Sorter100|5985_  = \new_Sorter100|5885_  & \new_Sorter100|5886_ ;
  assign \new_Sorter100|5986_  = \new_Sorter100|5885_  | \new_Sorter100|5886_ ;
  assign \new_Sorter100|5987_  = \new_Sorter100|5887_  & \new_Sorter100|5888_ ;
  assign \new_Sorter100|5988_  = \new_Sorter100|5887_  | \new_Sorter100|5888_ ;
  assign \new_Sorter100|5989_  = \new_Sorter100|5889_  & \new_Sorter100|5890_ ;
  assign \new_Sorter100|5990_  = \new_Sorter100|5889_  | \new_Sorter100|5890_ ;
  assign \new_Sorter100|5991_  = \new_Sorter100|5891_  & \new_Sorter100|5892_ ;
  assign \new_Sorter100|5992_  = \new_Sorter100|5891_  | \new_Sorter100|5892_ ;
  assign \new_Sorter100|5993_  = \new_Sorter100|5893_  & \new_Sorter100|5894_ ;
  assign \new_Sorter100|5994_  = \new_Sorter100|5893_  | \new_Sorter100|5894_ ;
  assign \new_Sorter100|5995_  = \new_Sorter100|5895_  & \new_Sorter100|5896_ ;
  assign \new_Sorter100|5996_  = \new_Sorter100|5895_  | \new_Sorter100|5896_ ;
  assign \new_Sorter100|5997_  = \new_Sorter100|5897_  & \new_Sorter100|5898_ ;
  assign \new_Sorter100|5998_  = \new_Sorter100|5897_  | \new_Sorter100|5898_ ;
  assign \new_Sorter100|6000_  = \new_Sorter100|5900_  & \new_Sorter100|5901_ ;
  assign \new_Sorter100|6001_  = \new_Sorter100|5900_  | \new_Sorter100|5901_ ;
  assign \new_Sorter100|6002_  = \new_Sorter100|5902_  & \new_Sorter100|5903_ ;
  assign \new_Sorter100|6003_  = \new_Sorter100|5902_  | \new_Sorter100|5903_ ;
  assign \new_Sorter100|6004_  = \new_Sorter100|5904_  & \new_Sorter100|5905_ ;
  assign \new_Sorter100|6005_  = \new_Sorter100|5904_  | \new_Sorter100|5905_ ;
  assign \new_Sorter100|6006_  = \new_Sorter100|5906_  & \new_Sorter100|5907_ ;
  assign \new_Sorter100|6007_  = \new_Sorter100|5906_  | \new_Sorter100|5907_ ;
  assign \new_Sorter100|6008_  = \new_Sorter100|5908_  & \new_Sorter100|5909_ ;
  assign \new_Sorter100|6009_  = \new_Sorter100|5908_  | \new_Sorter100|5909_ ;
  assign \new_Sorter100|6010_  = \new_Sorter100|5910_  & \new_Sorter100|5911_ ;
  assign \new_Sorter100|6011_  = \new_Sorter100|5910_  | \new_Sorter100|5911_ ;
  assign \new_Sorter100|6012_  = \new_Sorter100|5912_  & \new_Sorter100|5913_ ;
  assign \new_Sorter100|6013_  = \new_Sorter100|5912_  | \new_Sorter100|5913_ ;
  assign \new_Sorter100|6014_  = \new_Sorter100|5914_  & \new_Sorter100|5915_ ;
  assign \new_Sorter100|6015_  = \new_Sorter100|5914_  | \new_Sorter100|5915_ ;
  assign \new_Sorter100|6016_  = \new_Sorter100|5916_  & \new_Sorter100|5917_ ;
  assign \new_Sorter100|6017_  = \new_Sorter100|5916_  | \new_Sorter100|5917_ ;
  assign \new_Sorter100|6018_  = \new_Sorter100|5918_  & \new_Sorter100|5919_ ;
  assign \new_Sorter100|6019_  = \new_Sorter100|5918_  | \new_Sorter100|5919_ ;
  assign \new_Sorter100|6020_  = \new_Sorter100|5920_  & \new_Sorter100|5921_ ;
  assign \new_Sorter100|6021_  = \new_Sorter100|5920_  | \new_Sorter100|5921_ ;
  assign \new_Sorter100|6022_  = \new_Sorter100|5922_  & \new_Sorter100|5923_ ;
  assign \new_Sorter100|6023_  = \new_Sorter100|5922_  | \new_Sorter100|5923_ ;
  assign \new_Sorter100|6024_  = \new_Sorter100|5924_  & \new_Sorter100|5925_ ;
  assign \new_Sorter100|6025_  = \new_Sorter100|5924_  | \new_Sorter100|5925_ ;
  assign \new_Sorter100|6026_  = \new_Sorter100|5926_  & \new_Sorter100|5927_ ;
  assign \new_Sorter100|6027_  = \new_Sorter100|5926_  | \new_Sorter100|5927_ ;
  assign \new_Sorter100|6028_  = \new_Sorter100|5928_  & \new_Sorter100|5929_ ;
  assign \new_Sorter100|6029_  = \new_Sorter100|5928_  | \new_Sorter100|5929_ ;
  assign \new_Sorter100|6030_  = \new_Sorter100|5930_  & \new_Sorter100|5931_ ;
  assign \new_Sorter100|6031_  = \new_Sorter100|5930_  | \new_Sorter100|5931_ ;
  assign \new_Sorter100|6032_  = \new_Sorter100|5932_  & \new_Sorter100|5933_ ;
  assign \new_Sorter100|6033_  = \new_Sorter100|5932_  | \new_Sorter100|5933_ ;
  assign \new_Sorter100|6034_  = \new_Sorter100|5934_  & \new_Sorter100|5935_ ;
  assign \new_Sorter100|6035_  = \new_Sorter100|5934_  | \new_Sorter100|5935_ ;
  assign \new_Sorter100|6036_  = \new_Sorter100|5936_  & \new_Sorter100|5937_ ;
  assign \new_Sorter100|6037_  = \new_Sorter100|5936_  | \new_Sorter100|5937_ ;
  assign \new_Sorter100|6038_  = \new_Sorter100|5938_  & \new_Sorter100|5939_ ;
  assign \new_Sorter100|6039_  = \new_Sorter100|5938_  | \new_Sorter100|5939_ ;
  assign \new_Sorter100|6040_  = \new_Sorter100|5940_  & \new_Sorter100|5941_ ;
  assign \new_Sorter100|6041_  = \new_Sorter100|5940_  | \new_Sorter100|5941_ ;
  assign \new_Sorter100|6042_  = \new_Sorter100|5942_  & \new_Sorter100|5943_ ;
  assign \new_Sorter100|6043_  = \new_Sorter100|5942_  | \new_Sorter100|5943_ ;
  assign \new_Sorter100|6044_  = \new_Sorter100|5944_  & \new_Sorter100|5945_ ;
  assign \new_Sorter100|6045_  = \new_Sorter100|5944_  | \new_Sorter100|5945_ ;
  assign \new_Sorter100|6046_  = \new_Sorter100|5946_  & \new_Sorter100|5947_ ;
  assign \new_Sorter100|6047_  = \new_Sorter100|5946_  | \new_Sorter100|5947_ ;
  assign \new_Sorter100|6048_  = \new_Sorter100|5948_  & \new_Sorter100|5949_ ;
  assign \new_Sorter100|6049_  = \new_Sorter100|5948_  | \new_Sorter100|5949_ ;
  assign \new_Sorter100|6050_  = \new_Sorter100|5950_  & \new_Sorter100|5951_ ;
  assign \new_Sorter100|6051_  = \new_Sorter100|5950_  | \new_Sorter100|5951_ ;
  assign \new_Sorter100|6052_  = \new_Sorter100|5952_  & \new_Sorter100|5953_ ;
  assign \new_Sorter100|6053_  = \new_Sorter100|5952_  | \new_Sorter100|5953_ ;
  assign \new_Sorter100|6054_  = \new_Sorter100|5954_  & \new_Sorter100|5955_ ;
  assign \new_Sorter100|6055_  = \new_Sorter100|5954_  | \new_Sorter100|5955_ ;
  assign \new_Sorter100|6056_  = \new_Sorter100|5956_  & \new_Sorter100|5957_ ;
  assign \new_Sorter100|6057_  = \new_Sorter100|5956_  | \new_Sorter100|5957_ ;
  assign \new_Sorter100|6058_  = \new_Sorter100|5958_  & \new_Sorter100|5959_ ;
  assign \new_Sorter100|6059_  = \new_Sorter100|5958_  | \new_Sorter100|5959_ ;
  assign \new_Sorter100|6060_  = \new_Sorter100|5960_  & \new_Sorter100|5961_ ;
  assign \new_Sorter100|6061_  = \new_Sorter100|5960_  | \new_Sorter100|5961_ ;
  assign \new_Sorter100|6062_  = \new_Sorter100|5962_  & \new_Sorter100|5963_ ;
  assign \new_Sorter100|6063_  = \new_Sorter100|5962_  | \new_Sorter100|5963_ ;
  assign \new_Sorter100|6064_  = \new_Sorter100|5964_  & \new_Sorter100|5965_ ;
  assign \new_Sorter100|6065_  = \new_Sorter100|5964_  | \new_Sorter100|5965_ ;
  assign \new_Sorter100|6066_  = \new_Sorter100|5966_  & \new_Sorter100|5967_ ;
  assign \new_Sorter100|6067_  = \new_Sorter100|5966_  | \new_Sorter100|5967_ ;
  assign \new_Sorter100|6068_  = \new_Sorter100|5968_  & \new_Sorter100|5969_ ;
  assign \new_Sorter100|6069_  = \new_Sorter100|5968_  | \new_Sorter100|5969_ ;
  assign \new_Sorter100|6070_  = \new_Sorter100|5970_  & \new_Sorter100|5971_ ;
  assign \new_Sorter100|6071_  = \new_Sorter100|5970_  | \new_Sorter100|5971_ ;
  assign \new_Sorter100|6072_  = \new_Sorter100|5972_  & \new_Sorter100|5973_ ;
  assign \new_Sorter100|6073_  = \new_Sorter100|5972_  | \new_Sorter100|5973_ ;
  assign \new_Sorter100|6074_  = \new_Sorter100|5974_  & \new_Sorter100|5975_ ;
  assign \new_Sorter100|6075_  = \new_Sorter100|5974_  | \new_Sorter100|5975_ ;
  assign \new_Sorter100|6076_  = \new_Sorter100|5976_  & \new_Sorter100|5977_ ;
  assign \new_Sorter100|6077_  = \new_Sorter100|5976_  | \new_Sorter100|5977_ ;
  assign \new_Sorter100|6078_  = \new_Sorter100|5978_  & \new_Sorter100|5979_ ;
  assign \new_Sorter100|6079_  = \new_Sorter100|5978_  | \new_Sorter100|5979_ ;
  assign \new_Sorter100|6080_  = \new_Sorter100|5980_  & \new_Sorter100|5981_ ;
  assign \new_Sorter100|6081_  = \new_Sorter100|5980_  | \new_Sorter100|5981_ ;
  assign \new_Sorter100|6082_  = \new_Sorter100|5982_  & \new_Sorter100|5983_ ;
  assign \new_Sorter100|6083_  = \new_Sorter100|5982_  | \new_Sorter100|5983_ ;
  assign \new_Sorter100|6084_  = \new_Sorter100|5984_  & \new_Sorter100|5985_ ;
  assign \new_Sorter100|6085_  = \new_Sorter100|5984_  | \new_Sorter100|5985_ ;
  assign \new_Sorter100|6086_  = \new_Sorter100|5986_  & \new_Sorter100|5987_ ;
  assign \new_Sorter100|6087_  = \new_Sorter100|5986_  | \new_Sorter100|5987_ ;
  assign \new_Sorter100|6088_  = \new_Sorter100|5988_  & \new_Sorter100|5989_ ;
  assign \new_Sorter100|6089_  = \new_Sorter100|5988_  | \new_Sorter100|5989_ ;
  assign \new_Sorter100|6090_  = \new_Sorter100|5990_  & \new_Sorter100|5991_ ;
  assign \new_Sorter100|6091_  = \new_Sorter100|5990_  | \new_Sorter100|5991_ ;
  assign \new_Sorter100|6092_  = \new_Sorter100|5992_  & \new_Sorter100|5993_ ;
  assign \new_Sorter100|6093_  = \new_Sorter100|5992_  | \new_Sorter100|5993_ ;
  assign \new_Sorter100|6094_  = \new_Sorter100|5994_  & \new_Sorter100|5995_ ;
  assign \new_Sorter100|6095_  = \new_Sorter100|5994_  | \new_Sorter100|5995_ ;
  assign \new_Sorter100|6096_  = \new_Sorter100|5996_  & \new_Sorter100|5997_ ;
  assign \new_Sorter100|6097_  = \new_Sorter100|5996_  | \new_Sorter100|5997_ ;
  assign \new_Sorter100|6098_  = \new_Sorter100|5998_  & \new_Sorter100|5999_ ;
  assign \new_Sorter100|6099_  = \new_Sorter100|5998_  | \new_Sorter100|5999_ ;
  assign \new_Sorter100|6100_  = \new_Sorter100|6000_ ;
  assign \new_Sorter100|6199_  = \new_Sorter100|6099_ ;
  assign \new_Sorter100|6101_  = \new_Sorter100|6001_  & \new_Sorter100|6002_ ;
  assign \new_Sorter100|6102_  = \new_Sorter100|6001_  | \new_Sorter100|6002_ ;
  assign \new_Sorter100|6103_  = \new_Sorter100|6003_  & \new_Sorter100|6004_ ;
  assign \new_Sorter100|6104_  = \new_Sorter100|6003_  | \new_Sorter100|6004_ ;
  assign \new_Sorter100|6105_  = \new_Sorter100|6005_  & \new_Sorter100|6006_ ;
  assign \new_Sorter100|6106_  = \new_Sorter100|6005_  | \new_Sorter100|6006_ ;
  assign \new_Sorter100|6107_  = \new_Sorter100|6007_  & \new_Sorter100|6008_ ;
  assign \new_Sorter100|6108_  = \new_Sorter100|6007_  | \new_Sorter100|6008_ ;
  assign \new_Sorter100|6109_  = \new_Sorter100|6009_  & \new_Sorter100|6010_ ;
  assign \new_Sorter100|6110_  = \new_Sorter100|6009_  | \new_Sorter100|6010_ ;
  assign \new_Sorter100|6111_  = \new_Sorter100|6011_  & \new_Sorter100|6012_ ;
  assign \new_Sorter100|6112_  = \new_Sorter100|6011_  | \new_Sorter100|6012_ ;
  assign \new_Sorter100|6113_  = \new_Sorter100|6013_  & \new_Sorter100|6014_ ;
  assign \new_Sorter100|6114_  = \new_Sorter100|6013_  | \new_Sorter100|6014_ ;
  assign \new_Sorter100|6115_  = \new_Sorter100|6015_  & \new_Sorter100|6016_ ;
  assign \new_Sorter100|6116_  = \new_Sorter100|6015_  | \new_Sorter100|6016_ ;
  assign \new_Sorter100|6117_  = \new_Sorter100|6017_  & \new_Sorter100|6018_ ;
  assign \new_Sorter100|6118_  = \new_Sorter100|6017_  | \new_Sorter100|6018_ ;
  assign \new_Sorter100|6119_  = \new_Sorter100|6019_  & \new_Sorter100|6020_ ;
  assign \new_Sorter100|6120_  = \new_Sorter100|6019_  | \new_Sorter100|6020_ ;
  assign \new_Sorter100|6121_  = \new_Sorter100|6021_  & \new_Sorter100|6022_ ;
  assign \new_Sorter100|6122_  = \new_Sorter100|6021_  | \new_Sorter100|6022_ ;
  assign \new_Sorter100|6123_  = \new_Sorter100|6023_  & \new_Sorter100|6024_ ;
  assign \new_Sorter100|6124_  = \new_Sorter100|6023_  | \new_Sorter100|6024_ ;
  assign \new_Sorter100|6125_  = \new_Sorter100|6025_  & \new_Sorter100|6026_ ;
  assign \new_Sorter100|6126_  = \new_Sorter100|6025_  | \new_Sorter100|6026_ ;
  assign \new_Sorter100|6127_  = \new_Sorter100|6027_  & \new_Sorter100|6028_ ;
  assign \new_Sorter100|6128_  = \new_Sorter100|6027_  | \new_Sorter100|6028_ ;
  assign \new_Sorter100|6129_  = \new_Sorter100|6029_  & \new_Sorter100|6030_ ;
  assign \new_Sorter100|6130_  = \new_Sorter100|6029_  | \new_Sorter100|6030_ ;
  assign \new_Sorter100|6131_  = \new_Sorter100|6031_  & \new_Sorter100|6032_ ;
  assign \new_Sorter100|6132_  = \new_Sorter100|6031_  | \new_Sorter100|6032_ ;
  assign \new_Sorter100|6133_  = \new_Sorter100|6033_  & \new_Sorter100|6034_ ;
  assign \new_Sorter100|6134_  = \new_Sorter100|6033_  | \new_Sorter100|6034_ ;
  assign \new_Sorter100|6135_  = \new_Sorter100|6035_  & \new_Sorter100|6036_ ;
  assign \new_Sorter100|6136_  = \new_Sorter100|6035_  | \new_Sorter100|6036_ ;
  assign \new_Sorter100|6137_  = \new_Sorter100|6037_  & \new_Sorter100|6038_ ;
  assign \new_Sorter100|6138_  = \new_Sorter100|6037_  | \new_Sorter100|6038_ ;
  assign \new_Sorter100|6139_  = \new_Sorter100|6039_  & \new_Sorter100|6040_ ;
  assign \new_Sorter100|6140_  = \new_Sorter100|6039_  | \new_Sorter100|6040_ ;
  assign \new_Sorter100|6141_  = \new_Sorter100|6041_  & \new_Sorter100|6042_ ;
  assign \new_Sorter100|6142_  = \new_Sorter100|6041_  | \new_Sorter100|6042_ ;
  assign \new_Sorter100|6143_  = \new_Sorter100|6043_  & \new_Sorter100|6044_ ;
  assign \new_Sorter100|6144_  = \new_Sorter100|6043_  | \new_Sorter100|6044_ ;
  assign \new_Sorter100|6145_  = \new_Sorter100|6045_  & \new_Sorter100|6046_ ;
  assign \new_Sorter100|6146_  = \new_Sorter100|6045_  | \new_Sorter100|6046_ ;
  assign \new_Sorter100|6147_  = \new_Sorter100|6047_  & \new_Sorter100|6048_ ;
  assign \new_Sorter100|6148_  = \new_Sorter100|6047_  | \new_Sorter100|6048_ ;
  assign \new_Sorter100|6149_  = \new_Sorter100|6049_  & \new_Sorter100|6050_ ;
  assign \new_Sorter100|6150_  = \new_Sorter100|6049_  | \new_Sorter100|6050_ ;
  assign \new_Sorter100|6151_  = \new_Sorter100|6051_  & \new_Sorter100|6052_ ;
  assign \new_Sorter100|6152_  = \new_Sorter100|6051_  | \new_Sorter100|6052_ ;
  assign \new_Sorter100|6153_  = \new_Sorter100|6053_  & \new_Sorter100|6054_ ;
  assign \new_Sorter100|6154_  = \new_Sorter100|6053_  | \new_Sorter100|6054_ ;
  assign \new_Sorter100|6155_  = \new_Sorter100|6055_  & \new_Sorter100|6056_ ;
  assign \new_Sorter100|6156_  = \new_Sorter100|6055_  | \new_Sorter100|6056_ ;
  assign \new_Sorter100|6157_  = \new_Sorter100|6057_  & \new_Sorter100|6058_ ;
  assign \new_Sorter100|6158_  = \new_Sorter100|6057_  | \new_Sorter100|6058_ ;
  assign \new_Sorter100|6159_  = \new_Sorter100|6059_  & \new_Sorter100|6060_ ;
  assign \new_Sorter100|6160_  = \new_Sorter100|6059_  | \new_Sorter100|6060_ ;
  assign \new_Sorter100|6161_  = \new_Sorter100|6061_  & \new_Sorter100|6062_ ;
  assign \new_Sorter100|6162_  = \new_Sorter100|6061_  | \new_Sorter100|6062_ ;
  assign \new_Sorter100|6163_  = \new_Sorter100|6063_  & \new_Sorter100|6064_ ;
  assign \new_Sorter100|6164_  = \new_Sorter100|6063_  | \new_Sorter100|6064_ ;
  assign \new_Sorter100|6165_  = \new_Sorter100|6065_  & \new_Sorter100|6066_ ;
  assign \new_Sorter100|6166_  = \new_Sorter100|6065_  | \new_Sorter100|6066_ ;
  assign \new_Sorter100|6167_  = \new_Sorter100|6067_  & \new_Sorter100|6068_ ;
  assign \new_Sorter100|6168_  = \new_Sorter100|6067_  | \new_Sorter100|6068_ ;
  assign \new_Sorter100|6169_  = \new_Sorter100|6069_  & \new_Sorter100|6070_ ;
  assign \new_Sorter100|6170_  = \new_Sorter100|6069_  | \new_Sorter100|6070_ ;
  assign \new_Sorter100|6171_  = \new_Sorter100|6071_  & \new_Sorter100|6072_ ;
  assign \new_Sorter100|6172_  = \new_Sorter100|6071_  | \new_Sorter100|6072_ ;
  assign \new_Sorter100|6173_  = \new_Sorter100|6073_  & \new_Sorter100|6074_ ;
  assign \new_Sorter100|6174_  = \new_Sorter100|6073_  | \new_Sorter100|6074_ ;
  assign \new_Sorter100|6175_  = \new_Sorter100|6075_  & \new_Sorter100|6076_ ;
  assign \new_Sorter100|6176_  = \new_Sorter100|6075_  | \new_Sorter100|6076_ ;
  assign \new_Sorter100|6177_  = \new_Sorter100|6077_  & \new_Sorter100|6078_ ;
  assign \new_Sorter100|6178_  = \new_Sorter100|6077_  | \new_Sorter100|6078_ ;
  assign \new_Sorter100|6179_  = \new_Sorter100|6079_  & \new_Sorter100|6080_ ;
  assign \new_Sorter100|6180_  = \new_Sorter100|6079_  | \new_Sorter100|6080_ ;
  assign \new_Sorter100|6181_  = \new_Sorter100|6081_  & \new_Sorter100|6082_ ;
  assign \new_Sorter100|6182_  = \new_Sorter100|6081_  | \new_Sorter100|6082_ ;
  assign \new_Sorter100|6183_  = \new_Sorter100|6083_  & \new_Sorter100|6084_ ;
  assign \new_Sorter100|6184_  = \new_Sorter100|6083_  | \new_Sorter100|6084_ ;
  assign \new_Sorter100|6185_  = \new_Sorter100|6085_  & \new_Sorter100|6086_ ;
  assign \new_Sorter100|6186_  = \new_Sorter100|6085_  | \new_Sorter100|6086_ ;
  assign \new_Sorter100|6187_  = \new_Sorter100|6087_  & \new_Sorter100|6088_ ;
  assign \new_Sorter100|6188_  = \new_Sorter100|6087_  | \new_Sorter100|6088_ ;
  assign \new_Sorter100|6189_  = \new_Sorter100|6089_  & \new_Sorter100|6090_ ;
  assign \new_Sorter100|6190_  = \new_Sorter100|6089_  | \new_Sorter100|6090_ ;
  assign \new_Sorter100|6191_  = \new_Sorter100|6091_  & \new_Sorter100|6092_ ;
  assign \new_Sorter100|6192_  = \new_Sorter100|6091_  | \new_Sorter100|6092_ ;
  assign \new_Sorter100|6193_  = \new_Sorter100|6093_  & \new_Sorter100|6094_ ;
  assign \new_Sorter100|6194_  = \new_Sorter100|6093_  | \new_Sorter100|6094_ ;
  assign \new_Sorter100|6195_  = \new_Sorter100|6095_  & \new_Sorter100|6096_ ;
  assign \new_Sorter100|6196_  = \new_Sorter100|6095_  | \new_Sorter100|6096_ ;
  assign \new_Sorter100|6197_  = \new_Sorter100|6097_  & \new_Sorter100|6098_ ;
  assign \new_Sorter100|6198_  = \new_Sorter100|6097_  | \new_Sorter100|6098_ ;
  assign \new_Sorter100|6200_  = \new_Sorter100|6100_  & \new_Sorter100|6101_ ;
  assign \new_Sorter100|6201_  = \new_Sorter100|6100_  | \new_Sorter100|6101_ ;
  assign \new_Sorter100|6202_  = \new_Sorter100|6102_  & \new_Sorter100|6103_ ;
  assign \new_Sorter100|6203_  = \new_Sorter100|6102_  | \new_Sorter100|6103_ ;
  assign \new_Sorter100|6204_  = \new_Sorter100|6104_  & \new_Sorter100|6105_ ;
  assign \new_Sorter100|6205_  = \new_Sorter100|6104_  | \new_Sorter100|6105_ ;
  assign \new_Sorter100|6206_  = \new_Sorter100|6106_  & \new_Sorter100|6107_ ;
  assign \new_Sorter100|6207_  = \new_Sorter100|6106_  | \new_Sorter100|6107_ ;
  assign \new_Sorter100|6208_  = \new_Sorter100|6108_  & \new_Sorter100|6109_ ;
  assign \new_Sorter100|6209_  = \new_Sorter100|6108_  | \new_Sorter100|6109_ ;
  assign \new_Sorter100|6210_  = \new_Sorter100|6110_  & \new_Sorter100|6111_ ;
  assign \new_Sorter100|6211_  = \new_Sorter100|6110_  | \new_Sorter100|6111_ ;
  assign \new_Sorter100|6212_  = \new_Sorter100|6112_  & \new_Sorter100|6113_ ;
  assign \new_Sorter100|6213_  = \new_Sorter100|6112_  | \new_Sorter100|6113_ ;
  assign \new_Sorter100|6214_  = \new_Sorter100|6114_  & \new_Sorter100|6115_ ;
  assign \new_Sorter100|6215_  = \new_Sorter100|6114_  | \new_Sorter100|6115_ ;
  assign \new_Sorter100|6216_  = \new_Sorter100|6116_  & \new_Sorter100|6117_ ;
  assign \new_Sorter100|6217_  = \new_Sorter100|6116_  | \new_Sorter100|6117_ ;
  assign \new_Sorter100|6218_  = \new_Sorter100|6118_  & \new_Sorter100|6119_ ;
  assign \new_Sorter100|6219_  = \new_Sorter100|6118_  | \new_Sorter100|6119_ ;
  assign \new_Sorter100|6220_  = \new_Sorter100|6120_  & \new_Sorter100|6121_ ;
  assign \new_Sorter100|6221_  = \new_Sorter100|6120_  | \new_Sorter100|6121_ ;
  assign \new_Sorter100|6222_  = \new_Sorter100|6122_  & \new_Sorter100|6123_ ;
  assign \new_Sorter100|6223_  = \new_Sorter100|6122_  | \new_Sorter100|6123_ ;
  assign \new_Sorter100|6224_  = \new_Sorter100|6124_  & \new_Sorter100|6125_ ;
  assign \new_Sorter100|6225_  = \new_Sorter100|6124_  | \new_Sorter100|6125_ ;
  assign \new_Sorter100|6226_  = \new_Sorter100|6126_  & \new_Sorter100|6127_ ;
  assign \new_Sorter100|6227_  = \new_Sorter100|6126_  | \new_Sorter100|6127_ ;
  assign \new_Sorter100|6228_  = \new_Sorter100|6128_  & \new_Sorter100|6129_ ;
  assign \new_Sorter100|6229_  = \new_Sorter100|6128_  | \new_Sorter100|6129_ ;
  assign \new_Sorter100|6230_  = \new_Sorter100|6130_  & \new_Sorter100|6131_ ;
  assign \new_Sorter100|6231_  = \new_Sorter100|6130_  | \new_Sorter100|6131_ ;
  assign \new_Sorter100|6232_  = \new_Sorter100|6132_  & \new_Sorter100|6133_ ;
  assign \new_Sorter100|6233_  = \new_Sorter100|6132_  | \new_Sorter100|6133_ ;
  assign \new_Sorter100|6234_  = \new_Sorter100|6134_  & \new_Sorter100|6135_ ;
  assign \new_Sorter100|6235_  = \new_Sorter100|6134_  | \new_Sorter100|6135_ ;
  assign \new_Sorter100|6236_  = \new_Sorter100|6136_  & \new_Sorter100|6137_ ;
  assign \new_Sorter100|6237_  = \new_Sorter100|6136_  | \new_Sorter100|6137_ ;
  assign \new_Sorter100|6238_  = \new_Sorter100|6138_  & \new_Sorter100|6139_ ;
  assign \new_Sorter100|6239_  = \new_Sorter100|6138_  | \new_Sorter100|6139_ ;
  assign \new_Sorter100|6240_  = \new_Sorter100|6140_  & \new_Sorter100|6141_ ;
  assign \new_Sorter100|6241_  = \new_Sorter100|6140_  | \new_Sorter100|6141_ ;
  assign \new_Sorter100|6242_  = \new_Sorter100|6142_  & \new_Sorter100|6143_ ;
  assign \new_Sorter100|6243_  = \new_Sorter100|6142_  | \new_Sorter100|6143_ ;
  assign \new_Sorter100|6244_  = \new_Sorter100|6144_  & \new_Sorter100|6145_ ;
  assign \new_Sorter100|6245_  = \new_Sorter100|6144_  | \new_Sorter100|6145_ ;
  assign \new_Sorter100|6246_  = \new_Sorter100|6146_  & \new_Sorter100|6147_ ;
  assign \new_Sorter100|6247_  = \new_Sorter100|6146_  | \new_Sorter100|6147_ ;
  assign \new_Sorter100|6248_  = \new_Sorter100|6148_  & \new_Sorter100|6149_ ;
  assign \new_Sorter100|6249_  = \new_Sorter100|6148_  | \new_Sorter100|6149_ ;
  assign \new_Sorter100|6250_  = \new_Sorter100|6150_  & \new_Sorter100|6151_ ;
  assign \new_Sorter100|6251_  = \new_Sorter100|6150_  | \new_Sorter100|6151_ ;
  assign \new_Sorter100|6252_  = \new_Sorter100|6152_  & \new_Sorter100|6153_ ;
  assign \new_Sorter100|6253_  = \new_Sorter100|6152_  | \new_Sorter100|6153_ ;
  assign \new_Sorter100|6254_  = \new_Sorter100|6154_  & \new_Sorter100|6155_ ;
  assign \new_Sorter100|6255_  = \new_Sorter100|6154_  | \new_Sorter100|6155_ ;
  assign \new_Sorter100|6256_  = \new_Sorter100|6156_  & \new_Sorter100|6157_ ;
  assign \new_Sorter100|6257_  = \new_Sorter100|6156_  | \new_Sorter100|6157_ ;
  assign \new_Sorter100|6258_  = \new_Sorter100|6158_  & \new_Sorter100|6159_ ;
  assign \new_Sorter100|6259_  = \new_Sorter100|6158_  | \new_Sorter100|6159_ ;
  assign \new_Sorter100|6260_  = \new_Sorter100|6160_  & \new_Sorter100|6161_ ;
  assign \new_Sorter100|6261_  = \new_Sorter100|6160_  | \new_Sorter100|6161_ ;
  assign \new_Sorter100|6262_  = \new_Sorter100|6162_  & \new_Sorter100|6163_ ;
  assign \new_Sorter100|6263_  = \new_Sorter100|6162_  | \new_Sorter100|6163_ ;
  assign \new_Sorter100|6264_  = \new_Sorter100|6164_  & \new_Sorter100|6165_ ;
  assign \new_Sorter100|6265_  = \new_Sorter100|6164_  | \new_Sorter100|6165_ ;
  assign \new_Sorter100|6266_  = \new_Sorter100|6166_  & \new_Sorter100|6167_ ;
  assign \new_Sorter100|6267_  = \new_Sorter100|6166_  | \new_Sorter100|6167_ ;
  assign \new_Sorter100|6268_  = \new_Sorter100|6168_  & \new_Sorter100|6169_ ;
  assign \new_Sorter100|6269_  = \new_Sorter100|6168_  | \new_Sorter100|6169_ ;
  assign \new_Sorter100|6270_  = \new_Sorter100|6170_  & \new_Sorter100|6171_ ;
  assign \new_Sorter100|6271_  = \new_Sorter100|6170_  | \new_Sorter100|6171_ ;
  assign \new_Sorter100|6272_  = \new_Sorter100|6172_  & \new_Sorter100|6173_ ;
  assign \new_Sorter100|6273_  = \new_Sorter100|6172_  | \new_Sorter100|6173_ ;
  assign \new_Sorter100|6274_  = \new_Sorter100|6174_  & \new_Sorter100|6175_ ;
  assign \new_Sorter100|6275_  = \new_Sorter100|6174_  | \new_Sorter100|6175_ ;
  assign \new_Sorter100|6276_  = \new_Sorter100|6176_  & \new_Sorter100|6177_ ;
  assign \new_Sorter100|6277_  = \new_Sorter100|6176_  | \new_Sorter100|6177_ ;
  assign \new_Sorter100|6278_  = \new_Sorter100|6178_  & \new_Sorter100|6179_ ;
  assign \new_Sorter100|6279_  = \new_Sorter100|6178_  | \new_Sorter100|6179_ ;
  assign \new_Sorter100|6280_  = \new_Sorter100|6180_  & \new_Sorter100|6181_ ;
  assign \new_Sorter100|6281_  = \new_Sorter100|6180_  | \new_Sorter100|6181_ ;
  assign \new_Sorter100|6282_  = \new_Sorter100|6182_  & \new_Sorter100|6183_ ;
  assign \new_Sorter100|6283_  = \new_Sorter100|6182_  | \new_Sorter100|6183_ ;
  assign \new_Sorter100|6284_  = \new_Sorter100|6184_  & \new_Sorter100|6185_ ;
  assign \new_Sorter100|6285_  = \new_Sorter100|6184_  | \new_Sorter100|6185_ ;
  assign \new_Sorter100|6286_  = \new_Sorter100|6186_  & \new_Sorter100|6187_ ;
  assign \new_Sorter100|6287_  = \new_Sorter100|6186_  | \new_Sorter100|6187_ ;
  assign \new_Sorter100|6288_  = \new_Sorter100|6188_  & \new_Sorter100|6189_ ;
  assign \new_Sorter100|6289_  = \new_Sorter100|6188_  | \new_Sorter100|6189_ ;
  assign \new_Sorter100|6290_  = \new_Sorter100|6190_  & \new_Sorter100|6191_ ;
  assign \new_Sorter100|6291_  = \new_Sorter100|6190_  | \new_Sorter100|6191_ ;
  assign \new_Sorter100|6292_  = \new_Sorter100|6192_  & \new_Sorter100|6193_ ;
  assign \new_Sorter100|6293_  = \new_Sorter100|6192_  | \new_Sorter100|6193_ ;
  assign \new_Sorter100|6294_  = \new_Sorter100|6194_  & \new_Sorter100|6195_ ;
  assign \new_Sorter100|6295_  = \new_Sorter100|6194_  | \new_Sorter100|6195_ ;
  assign \new_Sorter100|6296_  = \new_Sorter100|6196_  & \new_Sorter100|6197_ ;
  assign \new_Sorter100|6297_  = \new_Sorter100|6196_  | \new_Sorter100|6197_ ;
  assign \new_Sorter100|6298_  = \new_Sorter100|6198_  & \new_Sorter100|6199_ ;
  assign \new_Sorter100|6299_  = \new_Sorter100|6198_  | \new_Sorter100|6199_ ;
  assign \new_Sorter100|6300_  = \new_Sorter100|6200_ ;
  assign \new_Sorter100|6399_  = \new_Sorter100|6299_ ;
  assign \new_Sorter100|6301_  = \new_Sorter100|6201_  & \new_Sorter100|6202_ ;
  assign \new_Sorter100|6302_  = \new_Sorter100|6201_  | \new_Sorter100|6202_ ;
  assign \new_Sorter100|6303_  = \new_Sorter100|6203_  & \new_Sorter100|6204_ ;
  assign \new_Sorter100|6304_  = \new_Sorter100|6203_  | \new_Sorter100|6204_ ;
  assign \new_Sorter100|6305_  = \new_Sorter100|6205_  & \new_Sorter100|6206_ ;
  assign \new_Sorter100|6306_  = \new_Sorter100|6205_  | \new_Sorter100|6206_ ;
  assign \new_Sorter100|6307_  = \new_Sorter100|6207_  & \new_Sorter100|6208_ ;
  assign \new_Sorter100|6308_  = \new_Sorter100|6207_  | \new_Sorter100|6208_ ;
  assign \new_Sorter100|6309_  = \new_Sorter100|6209_  & \new_Sorter100|6210_ ;
  assign \new_Sorter100|6310_  = \new_Sorter100|6209_  | \new_Sorter100|6210_ ;
  assign \new_Sorter100|6311_  = \new_Sorter100|6211_  & \new_Sorter100|6212_ ;
  assign \new_Sorter100|6312_  = \new_Sorter100|6211_  | \new_Sorter100|6212_ ;
  assign \new_Sorter100|6313_  = \new_Sorter100|6213_  & \new_Sorter100|6214_ ;
  assign \new_Sorter100|6314_  = \new_Sorter100|6213_  | \new_Sorter100|6214_ ;
  assign \new_Sorter100|6315_  = \new_Sorter100|6215_  & \new_Sorter100|6216_ ;
  assign \new_Sorter100|6316_  = \new_Sorter100|6215_  | \new_Sorter100|6216_ ;
  assign \new_Sorter100|6317_  = \new_Sorter100|6217_  & \new_Sorter100|6218_ ;
  assign \new_Sorter100|6318_  = \new_Sorter100|6217_  | \new_Sorter100|6218_ ;
  assign \new_Sorter100|6319_  = \new_Sorter100|6219_  & \new_Sorter100|6220_ ;
  assign \new_Sorter100|6320_  = \new_Sorter100|6219_  | \new_Sorter100|6220_ ;
  assign \new_Sorter100|6321_  = \new_Sorter100|6221_  & \new_Sorter100|6222_ ;
  assign \new_Sorter100|6322_  = \new_Sorter100|6221_  | \new_Sorter100|6222_ ;
  assign \new_Sorter100|6323_  = \new_Sorter100|6223_  & \new_Sorter100|6224_ ;
  assign \new_Sorter100|6324_  = \new_Sorter100|6223_  | \new_Sorter100|6224_ ;
  assign \new_Sorter100|6325_  = \new_Sorter100|6225_  & \new_Sorter100|6226_ ;
  assign \new_Sorter100|6326_  = \new_Sorter100|6225_  | \new_Sorter100|6226_ ;
  assign \new_Sorter100|6327_  = \new_Sorter100|6227_  & \new_Sorter100|6228_ ;
  assign \new_Sorter100|6328_  = \new_Sorter100|6227_  | \new_Sorter100|6228_ ;
  assign \new_Sorter100|6329_  = \new_Sorter100|6229_  & \new_Sorter100|6230_ ;
  assign \new_Sorter100|6330_  = \new_Sorter100|6229_  | \new_Sorter100|6230_ ;
  assign \new_Sorter100|6331_  = \new_Sorter100|6231_  & \new_Sorter100|6232_ ;
  assign \new_Sorter100|6332_  = \new_Sorter100|6231_  | \new_Sorter100|6232_ ;
  assign \new_Sorter100|6333_  = \new_Sorter100|6233_  & \new_Sorter100|6234_ ;
  assign \new_Sorter100|6334_  = \new_Sorter100|6233_  | \new_Sorter100|6234_ ;
  assign \new_Sorter100|6335_  = \new_Sorter100|6235_  & \new_Sorter100|6236_ ;
  assign \new_Sorter100|6336_  = \new_Sorter100|6235_  | \new_Sorter100|6236_ ;
  assign \new_Sorter100|6337_  = \new_Sorter100|6237_  & \new_Sorter100|6238_ ;
  assign \new_Sorter100|6338_  = \new_Sorter100|6237_  | \new_Sorter100|6238_ ;
  assign \new_Sorter100|6339_  = \new_Sorter100|6239_  & \new_Sorter100|6240_ ;
  assign \new_Sorter100|6340_  = \new_Sorter100|6239_  | \new_Sorter100|6240_ ;
  assign \new_Sorter100|6341_  = \new_Sorter100|6241_  & \new_Sorter100|6242_ ;
  assign \new_Sorter100|6342_  = \new_Sorter100|6241_  | \new_Sorter100|6242_ ;
  assign \new_Sorter100|6343_  = \new_Sorter100|6243_  & \new_Sorter100|6244_ ;
  assign \new_Sorter100|6344_  = \new_Sorter100|6243_  | \new_Sorter100|6244_ ;
  assign \new_Sorter100|6345_  = \new_Sorter100|6245_  & \new_Sorter100|6246_ ;
  assign \new_Sorter100|6346_  = \new_Sorter100|6245_  | \new_Sorter100|6246_ ;
  assign \new_Sorter100|6347_  = \new_Sorter100|6247_  & \new_Sorter100|6248_ ;
  assign \new_Sorter100|6348_  = \new_Sorter100|6247_  | \new_Sorter100|6248_ ;
  assign \new_Sorter100|6349_  = \new_Sorter100|6249_  & \new_Sorter100|6250_ ;
  assign \new_Sorter100|6350_  = \new_Sorter100|6249_  | \new_Sorter100|6250_ ;
  assign \new_Sorter100|6351_  = \new_Sorter100|6251_  & \new_Sorter100|6252_ ;
  assign \new_Sorter100|6352_  = \new_Sorter100|6251_  | \new_Sorter100|6252_ ;
  assign \new_Sorter100|6353_  = \new_Sorter100|6253_  & \new_Sorter100|6254_ ;
  assign \new_Sorter100|6354_  = \new_Sorter100|6253_  | \new_Sorter100|6254_ ;
  assign \new_Sorter100|6355_  = \new_Sorter100|6255_  & \new_Sorter100|6256_ ;
  assign \new_Sorter100|6356_  = \new_Sorter100|6255_  | \new_Sorter100|6256_ ;
  assign \new_Sorter100|6357_  = \new_Sorter100|6257_  & \new_Sorter100|6258_ ;
  assign \new_Sorter100|6358_  = \new_Sorter100|6257_  | \new_Sorter100|6258_ ;
  assign \new_Sorter100|6359_  = \new_Sorter100|6259_  & \new_Sorter100|6260_ ;
  assign \new_Sorter100|6360_  = \new_Sorter100|6259_  | \new_Sorter100|6260_ ;
  assign \new_Sorter100|6361_  = \new_Sorter100|6261_  & \new_Sorter100|6262_ ;
  assign \new_Sorter100|6362_  = \new_Sorter100|6261_  | \new_Sorter100|6262_ ;
  assign \new_Sorter100|6363_  = \new_Sorter100|6263_  & \new_Sorter100|6264_ ;
  assign \new_Sorter100|6364_  = \new_Sorter100|6263_  | \new_Sorter100|6264_ ;
  assign \new_Sorter100|6365_  = \new_Sorter100|6265_  & \new_Sorter100|6266_ ;
  assign \new_Sorter100|6366_  = \new_Sorter100|6265_  | \new_Sorter100|6266_ ;
  assign \new_Sorter100|6367_  = \new_Sorter100|6267_  & \new_Sorter100|6268_ ;
  assign \new_Sorter100|6368_  = \new_Sorter100|6267_  | \new_Sorter100|6268_ ;
  assign \new_Sorter100|6369_  = \new_Sorter100|6269_  & \new_Sorter100|6270_ ;
  assign \new_Sorter100|6370_  = \new_Sorter100|6269_  | \new_Sorter100|6270_ ;
  assign \new_Sorter100|6371_  = \new_Sorter100|6271_  & \new_Sorter100|6272_ ;
  assign \new_Sorter100|6372_  = \new_Sorter100|6271_  | \new_Sorter100|6272_ ;
  assign \new_Sorter100|6373_  = \new_Sorter100|6273_  & \new_Sorter100|6274_ ;
  assign \new_Sorter100|6374_  = \new_Sorter100|6273_  | \new_Sorter100|6274_ ;
  assign \new_Sorter100|6375_  = \new_Sorter100|6275_  & \new_Sorter100|6276_ ;
  assign \new_Sorter100|6376_  = \new_Sorter100|6275_  | \new_Sorter100|6276_ ;
  assign \new_Sorter100|6377_  = \new_Sorter100|6277_  & \new_Sorter100|6278_ ;
  assign \new_Sorter100|6378_  = \new_Sorter100|6277_  | \new_Sorter100|6278_ ;
  assign \new_Sorter100|6379_  = \new_Sorter100|6279_  & \new_Sorter100|6280_ ;
  assign \new_Sorter100|6380_  = \new_Sorter100|6279_  | \new_Sorter100|6280_ ;
  assign \new_Sorter100|6381_  = \new_Sorter100|6281_  & \new_Sorter100|6282_ ;
  assign \new_Sorter100|6382_  = \new_Sorter100|6281_  | \new_Sorter100|6282_ ;
  assign \new_Sorter100|6383_  = \new_Sorter100|6283_  & \new_Sorter100|6284_ ;
  assign \new_Sorter100|6384_  = \new_Sorter100|6283_  | \new_Sorter100|6284_ ;
  assign \new_Sorter100|6385_  = \new_Sorter100|6285_  & \new_Sorter100|6286_ ;
  assign \new_Sorter100|6386_  = \new_Sorter100|6285_  | \new_Sorter100|6286_ ;
  assign \new_Sorter100|6387_  = \new_Sorter100|6287_  & \new_Sorter100|6288_ ;
  assign \new_Sorter100|6388_  = \new_Sorter100|6287_  | \new_Sorter100|6288_ ;
  assign \new_Sorter100|6389_  = \new_Sorter100|6289_  & \new_Sorter100|6290_ ;
  assign \new_Sorter100|6390_  = \new_Sorter100|6289_  | \new_Sorter100|6290_ ;
  assign \new_Sorter100|6391_  = \new_Sorter100|6291_  & \new_Sorter100|6292_ ;
  assign \new_Sorter100|6392_  = \new_Sorter100|6291_  | \new_Sorter100|6292_ ;
  assign \new_Sorter100|6393_  = \new_Sorter100|6293_  & \new_Sorter100|6294_ ;
  assign \new_Sorter100|6394_  = \new_Sorter100|6293_  | \new_Sorter100|6294_ ;
  assign \new_Sorter100|6395_  = \new_Sorter100|6295_  & \new_Sorter100|6296_ ;
  assign \new_Sorter100|6396_  = \new_Sorter100|6295_  | \new_Sorter100|6296_ ;
  assign \new_Sorter100|6397_  = \new_Sorter100|6297_  & \new_Sorter100|6298_ ;
  assign \new_Sorter100|6398_  = \new_Sorter100|6297_  | \new_Sorter100|6298_ ;
  assign \new_Sorter100|6400_  = \new_Sorter100|6300_  & \new_Sorter100|6301_ ;
  assign \new_Sorter100|6401_  = \new_Sorter100|6300_  | \new_Sorter100|6301_ ;
  assign \new_Sorter100|6402_  = \new_Sorter100|6302_  & \new_Sorter100|6303_ ;
  assign \new_Sorter100|6403_  = \new_Sorter100|6302_  | \new_Sorter100|6303_ ;
  assign \new_Sorter100|6404_  = \new_Sorter100|6304_  & \new_Sorter100|6305_ ;
  assign \new_Sorter100|6405_  = \new_Sorter100|6304_  | \new_Sorter100|6305_ ;
  assign \new_Sorter100|6406_  = \new_Sorter100|6306_  & \new_Sorter100|6307_ ;
  assign \new_Sorter100|6407_  = \new_Sorter100|6306_  | \new_Sorter100|6307_ ;
  assign \new_Sorter100|6408_  = \new_Sorter100|6308_  & \new_Sorter100|6309_ ;
  assign \new_Sorter100|6409_  = \new_Sorter100|6308_  | \new_Sorter100|6309_ ;
  assign \new_Sorter100|6410_  = \new_Sorter100|6310_  & \new_Sorter100|6311_ ;
  assign \new_Sorter100|6411_  = \new_Sorter100|6310_  | \new_Sorter100|6311_ ;
  assign \new_Sorter100|6412_  = \new_Sorter100|6312_  & \new_Sorter100|6313_ ;
  assign \new_Sorter100|6413_  = \new_Sorter100|6312_  | \new_Sorter100|6313_ ;
  assign \new_Sorter100|6414_  = \new_Sorter100|6314_  & \new_Sorter100|6315_ ;
  assign \new_Sorter100|6415_  = \new_Sorter100|6314_  | \new_Sorter100|6315_ ;
  assign \new_Sorter100|6416_  = \new_Sorter100|6316_  & \new_Sorter100|6317_ ;
  assign \new_Sorter100|6417_  = \new_Sorter100|6316_  | \new_Sorter100|6317_ ;
  assign \new_Sorter100|6418_  = \new_Sorter100|6318_  & \new_Sorter100|6319_ ;
  assign \new_Sorter100|6419_  = \new_Sorter100|6318_  | \new_Sorter100|6319_ ;
  assign \new_Sorter100|6420_  = \new_Sorter100|6320_  & \new_Sorter100|6321_ ;
  assign \new_Sorter100|6421_  = \new_Sorter100|6320_  | \new_Sorter100|6321_ ;
  assign \new_Sorter100|6422_  = \new_Sorter100|6322_  & \new_Sorter100|6323_ ;
  assign \new_Sorter100|6423_  = \new_Sorter100|6322_  | \new_Sorter100|6323_ ;
  assign \new_Sorter100|6424_  = \new_Sorter100|6324_  & \new_Sorter100|6325_ ;
  assign \new_Sorter100|6425_  = \new_Sorter100|6324_  | \new_Sorter100|6325_ ;
  assign \new_Sorter100|6426_  = \new_Sorter100|6326_  & \new_Sorter100|6327_ ;
  assign \new_Sorter100|6427_  = \new_Sorter100|6326_  | \new_Sorter100|6327_ ;
  assign \new_Sorter100|6428_  = \new_Sorter100|6328_  & \new_Sorter100|6329_ ;
  assign \new_Sorter100|6429_  = \new_Sorter100|6328_  | \new_Sorter100|6329_ ;
  assign \new_Sorter100|6430_  = \new_Sorter100|6330_  & \new_Sorter100|6331_ ;
  assign \new_Sorter100|6431_  = \new_Sorter100|6330_  | \new_Sorter100|6331_ ;
  assign \new_Sorter100|6432_  = \new_Sorter100|6332_  & \new_Sorter100|6333_ ;
  assign \new_Sorter100|6433_  = \new_Sorter100|6332_  | \new_Sorter100|6333_ ;
  assign \new_Sorter100|6434_  = \new_Sorter100|6334_  & \new_Sorter100|6335_ ;
  assign \new_Sorter100|6435_  = \new_Sorter100|6334_  | \new_Sorter100|6335_ ;
  assign \new_Sorter100|6436_  = \new_Sorter100|6336_  & \new_Sorter100|6337_ ;
  assign \new_Sorter100|6437_  = \new_Sorter100|6336_  | \new_Sorter100|6337_ ;
  assign \new_Sorter100|6438_  = \new_Sorter100|6338_  & \new_Sorter100|6339_ ;
  assign \new_Sorter100|6439_  = \new_Sorter100|6338_  | \new_Sorter100|6339_ ;
  assign \new_Sorter100|6440_  = \new_Sorter100|6340_  & \new_Sorter100|6341_ ;
  assign \new_Sorter100|6441_  = \new_Sorter100|6340_  | \new_Sorter100|6341_ ;
  assign \new_Sorter100|6442_  = \new_Sorter100|6342_  & \new_Sorter100|6343_ ;
  assign \new_Sorter100|6443_  = \new_Sorter100|6342_  | \new_Sorter100|6343_ ;
  assign \new_Sorter100|6444_  = \new_Sorter100|6344_  & \new_Sorter100|6345_ ;
  assign \new_Sorter100|6445_  = \new_Sorter100|6344_  | \new_Sorter100|6345_ ;
  assign \new_Sorter100|6446_  = \new_Sorter100|6346_  & \new_Sorter100|6347_ ;
  assign \new_Sorter100|6447_  = \new_Sorter100|6346_  | \new_Sorter100|6347_ ;
  assign \new_Sorter100|6448_  = \new_Sorter100|6348_  & \new_Sorter100|6349_ ;
  assign \new_Sorter100|6449_  = \new_Sorter100|6348_  | \new_Sorter100|6349_ ;
  assign \new_Sorter100|6450_  = \new_Sorter100|6350_  & \new_Sorter100|6351_ ;
  assign \new_Sorter100|6451_  = \new_Sorter100|6350_  | \new_Sorter100|6351_ ;
  assign \new_Sorter100|6452_  = \new_Sorter100|6352_  & \new_Sorter100|6353_ ;
  assign \new_Sorter100|6453_  = \new_Sorter100|6352_  | \new_Sorter100|6353_ ;
  assign \new_Sorter100|6454_  = \new_Sorter100|6354_  & \new_Sorter100|6355_ ;
  assign \new_Sorter100|6455_  = \new_Sorter100|6354_  | \new_Sorter100|6355_ ;
  assign \new_Sorter100|6456_  = \new_Sorter100|6356_  & \new_Sorter100|6357_ ;
  assign \new_Sorter100|6457_  = \new_Sorter100|6356_  | \new_Sorter100|6357_ ;
  assign \new_Sorter100|6458_  = \new_Sorter100|6358_  & \new_Sorter100|6359_ ;
  assign \new_Sorter100|6459_  = \new_Sorter100|6358_  | \new_Sorter100|6359_ ;
  assign \new_Sorter100|6460_  = \new_Sorter100|6360_  & \new_Sorter100|6361_ ;
  assign \new_Sorter100|6461_  = \new_Sorter100|6360_  | \new_Sorter100|6361_ ;
  assign \new_Sorter100|6462_  = \new_Sorter100|6362_  & \new_Sorter100|6363_ ;
  assign \new_Sorter100|6463_  = \new_Sorter100|6362_  | \new_Sorter100|6363_ ;
  assign \new_Sorter100|6464_  = \new_Sorter100|6364_  & \new_Sorter100|6365_ ;
  assign \new_Sorter100|6465_  = \new_Sorter100|6364_  | \new_Sorter100|6365_ ;
  assign \new_Sorter100|6466_  = \new_Sorter100|6366_  & \new_Sorter100|6367_ ;
  assign \new_Sorter100|6467_  = \new_Sorter100|6366_  | \new_Sorter100|6367_ ;
  assign \new_Sorter100|6468_  = \new_Sorter100|6368_  & \new_Sorter100|6369_ ;
  assign \new_Sorter100|6469_  = \new_Sorter100|6368_  | \new_Sorter100|6369_ ;
  assign \new_Sorter100|6470_  = \new_Sorter100|6370_  & \new_Sorter100|6371_ ;
  assign \new_Sorter100|6471_  = \new_Sorter100|6370_  | \new_Sorter100|6371_ ;
  assign \new_Sorter100|6472_  = \new_Sorter100|6372_  & \new_Sorter100|6373_ ;
  assign \new_Sorter100|6473_  = \new_Sorter100|6372_  | \new_Sorter100|6373_ ;
  assign \new_Sorter100|6474_  = \new_Sorter100|6374_  & \new_Sorter100|6375_ ;
  assign \new_Sorter100|6475_  = \new_Sorter100|6374_  | \new_Sorter100|6375_ ;
  assign \new_Sorter100|6476_  = \new_Sorter100|6376_  & \new_Sorter100|6377_ ;
  assign \new_Sorter100|6477_  = \new_Sorter100|6376_  | \new_Sorter100|6377_ ;
  assign \new_Sorter100|6478_  = \new_Sorter100|6378_  & \new_Sorter100|6379_ ;
  assign \new_Sorter100|6479_  = \new_Sorter100|6378_  | \new_Sorter100|6379_ ;
  assign \new_Sorter100|6480_  = \new_Sorter100|6380_  & \new_Sorter100|6381_ ;
  assign \new_Sorter100|6481_  = \new_Sorter100|6380_  | \new_Sorter100|6381_ ;
  assign \new_Sorter100|6482_  = \new_Sorter100|6382_  & \new_Sorter100|6383_ ;
  assign \new_Sorter100|6483_  = \new_Sorter100|6382_  | \new_Sorter100|6383_ ;
  assign \new_Sorter100|6484_  = \new_Sorter100|6384_  & \new_Sorter100|6385_ ;
  assign \new_Sorter100|6485_  = \new_Sorter100|6384_  | \new_Sorter100|6385_ ;
  assign \new_Sorter100|6486_  = \new_Sorter100|6386_  & \new_Sorter100|6387_ ;
  assign \new_Sorter100|6487_  = \new_Sorter100|6386_  | \new_Sorter100|6387_ ;
  assign \new_Sorter100|6488_  = \new_Sorter100|6388_  & \new_Sorter100|6389_ ;
  assign \new_Sorter100|6489_  = \new_Sorter100|6388_  | \new_Sorter100|6389_ ;
  assign \new_Sorter100|6490_  = \new_Sorter100|6390_  & \new_Sorter100|6391_ ;
  assign \new_Sorter100|6491_  = \new_Sorter100|6390_  | \new_Sorter100|6391_ ;
  assign \new_Sorter100|6492_  = \new_Sorter100|6392_  & \new_Sorter100|6393_ ;
  assign \new_Sorter100|6493_  = \new_Sorter100|6392_  | \new_Sorter100|6393_ ;
  assign \new_Sorter100|6494_  = \new_Sorter100|6394_  & \new_Sorter100|6395_ ;
  assign \new_Sorter100|6495_  = \new_Sorter100|6394_  | \new_Sorter100|6395_ ;
  assign \new_Sorter100|6496_  = \new_Sorter100|6396_  & \new_Sorter100|6397_ ;
  assign \new_Sorter100|6497_  = \new_Sorter100|6396_  | \new_Sorter100|6397_ ;
  assign \new_Sorter100|6498_  = \new_Sorter100|6398_  & \new_Sorter100|6399_ ;
  assign \new_Sorter100|6499_  = \new_Sorter100|6398_  | \new_Sorter100|6399_ ;
  assign \new_Sorter100|6500_  = \new_Sorter100|6400_ ;
  assign \new_Sorter100|6599_  = \new_Sorter100|6499_ ;
  assign \new_Sorter100|6501_  = \new_Sorter100|6401_  & \new_Sorter100|6402_ ;
  assign \new_Sorter100|6502_  = \new_Sorter100|6401_  | \new_Sorter100|6402_ ;
  assign \new_Sorter100|6503_  = \new_Sorter100|6403_  & \new_Sorter100|6404_ ;
  assign \new_Sorter100|6504_  = \new_Sorter100|6403_  | \new_Sorter100|6404_ ;
  assign \new_Sorter100|6505_  = \new_Sorter100|6405_  & \new_Sorter100|6406_ ;
  assign \new_Sorter100|6506_  = \new_Sorter100|6405_  | \new_Sorter100|6406_ ;
  assign \new_Sorter100|6507_  = \new_Sorter100|6407_  & \new_Sorter100|6408_ ;
  assign \new_Sorter100|6508_  = \new_Sorter100|6407_  | \new_Sorter100|6408_ ;
  assign \new_Sorter100|6509_  = \new_Sorter100|6409_  & \new_Sorter100|6410_ ;
  assign \new_Sorter100|6510_  = \new_Sorter100|6409_  | \new_Sorter100|6410_ ;
  assign \new_Sorter100|6511_  = \new_Sorter100|6411_  & \new_Sorter100|6412_ ;
  assign \new_Sorter100|6512_  = \new_Sorter100|6411_  | \new_Sorter100|6412_ ;
  assign \new_Sorter100|6513_  = \new_Sorter100|6413_  & \new_Sorter100|6414_ ;
  assign \new_Sorter100|6514_  = \new_Sorter100|6413_  | \new_Sorter100|6414_ ;
  assign \new_Sorter100|6515_  = \new_Sorter100|6415_  & \new_Sorter100|6416_ ;
  assign \new_Sorter100|6516_  = \new_Sorter100|6415_  | \new_Sorter100|6416_ ;
  assign \new_Sorter100|6517_  = \new_Sorter100|6417_  & \new_Sorter100|6418_ ;
  assign \new_Sorter100|6518_  = \new_Sorter100|6417_  | \new_Sorter100|6418_ ;
  assign \new_Sorter100|6519_  = \new_Sorter100|6419_  & \new_Sorter100|6420_ ;
  assign \new_Sorter100|6520_  = \new_Sorter100|6419_  | \new_Sorter100|6420_ ;
  assign \new_Sorter100|6521_  = \new_Sorter100|6421_  & \new_Sorter100|6422_ ;
  assign \new_Sorter100|6522_  = \new_Sorter100|6421_  | \new_Sorter100|6422_ ;
  assign \new_Sorter100|6523_  = \new_Sorter100|6423_  & \new_Sorter100|6424_ ;
  assign \new_Sorter100|6524_  = \new_Sorter100|6423_  | \new_Sorter100|6424_ ;
  assign \new_Sorter100|6525_  = \new_Sorter100|6425_  & \new_Sorter100|6426_ ;
  assign \new_Sorter100|6526_  = \new_Sorter100|6425_  | \new_Sorter100|6426_ ;
  assign \new_Sorter100|6527_  = \new_Sorter100|6427_  & \new_Sorter100|6428_ ;
  assign \new_Sorter100|6528_  = \new_Sorter100|6427_  | \new_Sorter100|6428_ ;
  assign \new_Sorter100|6529_  = \new_Sorter100|6429_  & \new_Sorter100|6430_ ;
  assign \new_Sorter100|6530_  = \new_Sorter100|6429_  | \new_Sorter100|6430_ ;
  assign \new_Sorter100|6531_  = \new_Sorter100|6431_  & \new_Sorter100|6432_ ;
  assign \new_Sorter100|6532_  = \new_Sorter100|6431_  | \new_Sorter100|6432_ ;
  assign \new_Sorter100|6533_  = \new_Sorter100|6433_  & \new_Sorter100|6434_ ;
  assign \new_Sorter100|6534_  = \new_Sorter100|6433_  | \new_Sorter100|6434_ ;
  assign \new_Sorter100|6535_  = \new_Sorter100|6435_  & \new_Sorter100|6436_ ;
  assign \new_Sorter100|6536_  = \new_Sorter100|6435_  | \new_Sorter100|6436_ ;
  assign \new_Sorter100|6537_  = \new_Sorter100|6437_  & \new_Sorter100|6438_ ;
  assign \new_Sorter100|6538_  = \new_Sorter100|6437_  | \new_Sorter100|6438_ ;
  assign \new_Sorter100|6539_  = \new_Sorter100|6439_  & \new_Sorter100|6440_ ;
  assign \new_Sorter100|6540_  = \new_Sorter100|6439_  | \new_Sorter100|6440_ ;
  assign \new_Sorter100|6541_  = \new_Sorter100|6441_  & \new_Sorter100|6442_ ;
  assign \new_Sorter100|6542_  = \new_Sorter100|6441_  | \new_Sorter100|6442_ ;
  assign \new_Sorter100|6543_  = \new_Sorter100|6443_  & \new_Sorter100|6444_ ;
  assign \new_Sorter100|6544_  = \new_Sorter100|6443_  | \new_Sorter100|6444_ ;
  assign \new_Sorter100|6545_  = \new_Sorter100|6445_  & \new_Sorter100|6446_ ;
  assign \new_Sorter100|6546_  = \new_Sorter100|6445_  | \new_Sorter100|6446_ ;
  assign \new_Sorter100|6547_  = \new_Sorter100|6447_  & \new_Sorter100|6448_ ;
  assign \new_Sorter100|6548_  = \new_Sorter100|6447_  | \new_Sorter100|6448_ ;
  assign \new_Sorter100|6549_  = \new_Sorter100|6449_  & \new_Sorter100|6450_ ;
  assign \new_Sorter100|6550_  = \new_Sorter100|6449_  | \new_Sorter100|6450_ ;
  assign \new_Sorter100|6551_  = \new_Sorter100|6451_  & \new_Sorter100|6452_ ;
  assign \new_Sorter100|6552_  = \new_Sorter100|6451_  | \new_Sorter100|6452_ ;
  assign \new_Sorter100|6553_  = \new_Sorter100|6453_  & \new_Sorter100|6454_ ;
  assign \new_Sorter100|6554_  = \new_Sorter100|6453_  | \new_Sorter100|6454_ ;
  assign \new_Sorter100|6555_  = \new_Sorter100|6455_  & \new_Sorter100|6456_ ;
  assign \new_Sorter100|6556_  = \new_Sorter100|6455_  | \new_Sorter100|6456_ ;
  assign \new_Sorter100|6557_  = \new_Sorter100|6457_  & \new_Sorter100|6458_ ;
  assign \new_Sorter100|6558_  = \new_Sorter100|6457_  | \new_Sorter100|6458_ ;
  assign \new_Sorter100|6559_  = \new_Sorter100|6459_  & \new_Sorter100|6460_ ;
  assign \new_Sorter100|6560_  = \new_Sorter100|6459_  | \new_Sorter100|6460_ ;
  assign \new_Sorter100|6561_  = \new_Sorter100|6461_  & \new_Sorter100|6462_ ;
  assign \new_Sorter100|6562_  = \new_Sorter100|6461_  | \new_Sorter100|6462_ ;
  assign \new_Sorter100|6563_  = \new_Sorter100|6463_  & \new_Sorter100|6464_ ;
  assign \new_Sorter100|6564_  = \new_Sorter100|6463_  | \new_Sorter100|6464_ ;
  assign \new_Sorter100|6565_  = \new_Sorter100|6465_  & \new_Sorter100|6466_ ;
  assign \new_Sorter100|6566_  = \new_Sorter100|6465_  | \new_Sorter100|6466_ ;
  assign \new_Sorter100|6567_  = \new_Sorter100|6467_  & \new_Sorter100|6468_ ;
  assign \new_Sorter100|6568_  = \new_Sorter100|6467_  | \new_Sorter100|6468_ ;
  assign \new_Sorter100|6569_  = \new_Sorter100|6469_  & \new_Sorter100|6470_ ;
  assign \new_Sorter100|6570_  = \new_Sorter100|6469_  | \new_Sorter100|6470_ ;
  assign \new_Sorter100|6571_  = \new_Sorter100|6471_  & \new_Sorter100|6472_ ;
  assign \new_Sorter100|6572_  = \new_Sorter100|6471_  | \new_Sorter100|6472_ ;
  assign \new_Sorter100|6573_  = \new_Sorter100|6473_  & \new_Sorter100|6474_ ;
  assign \new_Sorter100|6574_  = \new_Sorter100|6473_  | \new_Sorter100|6474_ ;
  assign \new_Sorter100|6575_  = \new_Sorter100|6475_  & \new_Sorter100|6476_ ;
  assign \new_Sorter100|6576_  = \new_Sorter100|6475_  | \new_Sorter100|6476_ ;
  assign \new_Sorter100|6577_  = \new_Sorter100|6477_  & \new_Sorter100|6478_ ;
  assign \new_Sorter100|6578_  = \new_Sorter100|6477_  | \new_Sorter100|6478_ ;
  assign \new_Sorter100|6579_  = \new_Sorter100|6479_  & \new_Sorter100|6480_ ;
  assign \new_Sorter100|6580_  = \new_Sorter100|6479_  | \new_Sorter100|6480_ ;
  assign \new_Sorter100|6581_  = \new_Sorter100|6481_  & \new_Sorter100|6482_ ;
  assign \new_Sorter100|6582_  = \new_Sorter100|6481_  | \new_Sorter100|6482_ ;
  assign \new_Sorter100|6583_  = \new_Sorter100|6483_  & \new_Sorter100|6484_ ;
  assign \new_Sorter100|6584_  = \new_Sorter100|6483_  | \new_Sorter100|6484_ ;
  assign \new_Sorter100|6585_  = \new_Sorter100|6485_  & \new_Sorter100|6486_ ;
  assign \new_Sorter100|6586_  = \new_Sorter100|6485_  | \new_Sorter100|6486_ ;
  assign \new_Sorter100|6587_  = \new_Sorter100|6487_  & \new_Sorter100|6488_ ;
  assign \new_Sorter100|6588_  = \new_Sorter100|6487_  | \new_Sorter100|6488_ ;
  assign \new_Sorter100|6589_  = \new_Sorter100|6489_  & \new_Sorter100|6490_ ;
  assign \new_Sorter100|6590_  = \new_Sorter100|6489_  | \new_Sorter100|6490_ ;
  assign \new_Sorter100|6591_  = \new_Sorter100|6491_  & \new_Sorter100|6492_ ;
  assign \new_Sorter100|6592_  = \new_Sorter100|6491_  | \new_Sorter100|6492_ ;
  assign \new_Sorter100|6593_  = \new_Sorter100|6493_  & \new_Sorter100|6494_ ;
  assign \new_Sorter100|6594_  = \new_Sorter100|6493_  | \new_Sorter100|6494_ ;
  assign \new_Sorter100|6595_  = \new_Sorter100|6495_  & \new_Sorter100|6496_ ;
  assign \new_Sorter100|6596_  = \new_Sorter100|6495_  | \new_Sorter100|6496_ ;
  assign \new_Sorter100|6597_  = \new_Sorter100|6497_  & \new_Sorter100|6498_ ;
  assign \new_Sorter100|6598_  = \new_Sorter100|6497_  | \new_Sorter100|6498_ ;
  assign \new_Sorter100|6600_  = \new_Sorter100|6500_  & \new_Sorter100|6501_ ;
  assign \new_Sorter100|6601_  = \new_Sorter100|6500_  | \new_Sorter100|6501_ ;
  assign \new_Sorter100|6602_  = \new_Sorter100|6502_  & \new_Sorter100|6503_ ;
  assign \new_Sorter100|6603_  = \new_Sorter100|6502_  | \new_Sorter100|6503_ ;
  assign \new_Sorter100|6604_  = \new_Sorter100|6504_  & \new_Sorter100|6505_ ;
  assign \new_Sorter100|6605_  = \new_Sorter100|6504_  | \new_Sorter100|6505_ ;
  assign \new_Sorter100|6606_  = \new_Sorter100|6506_  & \new_Sorter100|6507_ ;
  assign \new_Sorter100|6607_  = \new_Sorter100|6506_  | \new_Sorter100|6507_ ;
  assign \new_Sorter100|6608_  = \new_Sorter100|6508_  & \new_Sorter100|6509_ ;
  assign \new_Sorter100|6609_  = \new_Sorter100|6508_  | \new_Sorter100|6509_ ;
  assign \new_Sorter100|6610_  = \new_Sorter100|6510_  & \new_Sorter100|6511_ ;
  assign \new_Sorter100|6611_  = \new_Sorter100|6510_  | \new_Sorter100|6511_ ;
  assign \new_Sorter100|6612_  = \new_Sorter100|6512_  & \new_Sorter100|6513_ ;
  assign \new_Sorter100|6613_  = \new_Sorter100|6512_  | \new_Sorter100|6513_ ;
  assign \new_Sorter100|6614_  = \new_Sorter100|6514_  & \new_Sorter100|6515_ ;
  assign \new_Sorter100|6615_  = \new_Sorter100|6514_  | \new_Sorter100|6515_ ;
  assign \new_Sorter100|6616_  = \new_Sorter100|6516_  & \new_Sorter100|6517_ ;
  assign \new_Sorter100|6617_  = \new_Sorter100|6516_  | \new_Sorter100|6517_ ;
  assign \new_Sorter100|6618_  = \new_Sorter100|6518_  & \new_Sorter100|6519_ ;
  assign \new_Sorter100|6619_  = \new_Sorter100|6518_  | \new_Sorter100|6519_ ;
  assign \new_Sorter100|6620_  = \new_Sorter100|6520_  & \new_Sorter100|6521_ ;
  assign \new_Sorter100|6621_  = \new_Sorter100|6520_  | \new_Sorter100|6521_ ;
  assign \new_Sorter100|6622_  = \new_Sorter100|6522_  & \new_Sorter100|6523_ ;
  assign \new_Sorter100|6623_  = \new_Sorter100|6522_  | \new_Sorter100|6523_ ;
  assign \new_Sorter100|6624_  = \new_Sorter100|6524_  & \new_Sorter100|6525_ ;
  assign \new_Sorter100|6625_  = \new_Sorter100|6524_  | \new_Sorter100|6525_ ;
  assign \new_Sorter100|6626_  = \new_Sorter100|6526_  & \new_Sorter100|6527_ ;
  assign \new_Sorter100|6627_  = \new_Sorter100|6526_  | \new_Sorter100|6527_ ;
  assign \new_Sorter100|6628_  = \new_Sorter100|6528_  & \new_Sorter100|6529_ ;
  assign \new_Sorter100|6629_  = \new_Sorter100|6528_  | \new_Sorter100|6529_ ;
  assign \new_Sorter100|6630_  = \new_Sorter100|6530_  & \new_Sorter100|6531_ ;
  assign \new_Sorter100|6631_  = \new_Sorter100|6530_  | \new_Sorter100|6531_ ;
  assign \new_Sorter100|6632_  = \new_Sorter100|6532_  & \new_Sorter100|6533_ ;
  assign \new_Sorter100|6633_  = \new_Sorter100|6532_  | \new_Sorter100|6533_ ;
  assign \new_Sorter100|6634_  = \new_Sorter100|6534_  & \new_Sorter100|6535_ ;
  assign \new_Sorter100|6635_  = \new_Sorter100|6534_  | \new_Sorter100|6535_ ;
  assign \new_Sorter100|6636_  = \new_Sorter100|6536_  & \new_Sorter100|6537_ ;
  assign \new_Sorter100|6637_  = \new_Sorter100|6536_  | \new_Sorter100|6537_ ;
  assign \new_Sorter100|6638_  = \new_Sorter100|6538_  & \new_Sorter100|6539_ ;
  assign \new_Sorter100|6639_  = \new_Sorter100|6538_  | \new_Sorter100|6539_ ;
  assign \new_Sorter100|6640_  = \new_Sorter100|6540_  & \new_Sorter100|6541_ ;
  assign \new_Sorter100|6641_  = \new_Sorter100|6540_  | \new_Sorter100|6541_ ;
  assign \new_Sorter100|6642_  = \new_Sorter100|6542_  & \new_Sorter100|6543_ ;
  assign \new_Sorter100|6643_  = \new_Sorter100|6542_  | \new_Sorter100|6543_ ;
  assign \new_Sorter100|6644_  = \new_Sorter100|6544_  & \new_Sorter100|6545_ ;
  assign \new_Sorter100|6645_  = \new_Sorter100|6544_  | \new_Sorter100|6545_ ;
  assign \new_Sorter100|6646_  = \new_Sorter100|6546_  & \new_Sorter100|6547_ ;
  assign \new_Sorter100|6647_  = \new_Sorter100|6546_  | \new_Sorter100|6547_ ;
  assign \new_Sorter100|6648_  = \new_Sorter100|6548_  & \new_Sorter100|6549_ ;
  assign \new_Sorter100|6649_  = \new_Sorter100|6548_  | \new_Sorter100|6549_ ;
  assign \new_Sorter100|6650_  = \new_Sorter100|6550_  & \new_Sorter100|6551_ ;
  assign \new_Sorter100|6651_  = \new_Sorter100|6550_  | \new_Sorter100|6551_ ;
  assign \new_Sorter100|6652_  = \new_Sorter100|6552_  & \new_Sorter100|6553_ ;
  assign \new_Sorter100|6653_  = \new_Sorter100|6552_  | \new_Sorter100|6553_ ;
  assign \new_Sorter100|6654_  = \new_Sorter100|6554_  & \new_Sorter100|6555_ ;
  assign \new_Sorter100|6655_  = \new_Sorter100|6554_  | \new_Sorter100|6555_ ;
  assign \new_Sorter100|6656_  = \new_Sorter100|6556_  & \new_Sorter100|6557_ ;
  assign \new_Sorter100|6657_  = \new_Sorter100|6556_  | \new_Sorter100|6557_ ;
  assign \new_Sorter100|6658_  = \new_Sorter100|6558_  & \new_Sorter100|6559_ ;
  assign \new_Sorter100|6659_  = \new_Sorter100|6558_  | \new_Sorter100|6559_ ;
  assign \new_Sorter100|6660_  = \new_Sorter100|6560_  & \new_Sorter100|6561_ ;
  assign \new_Sorter100|6661_  = \new_Sorter100|6560_  | \new_Sorter100|6561_ ;
  assign \new_Sorter100|6662_  = \new_Sorter100|6562_  & \new_Sorter100|6563_ ;
  assign \new_Sorter100|6663_  = \new_Sorter100|6562_  | \new_Sorter100|6563_ ;
  assign \new_Sorter100|6664_  = \new_Sorter100|6564_  & \new_Sorter100|6565_ ;
  assign \new_Sorter100|6665_  = \new_Sorter100|6564_  | \new_Sorter100|6565_ ;
  assign \new_Sorter100|6666_  = \new_Sorter100|6566_  & \new_Sorter100|6567_ ;
  assign \new_Sorter100|6667_  = \new_Sorter100|6566_  | \new_Sorter100|6567_ ;
  assign \new_Sorter100|6668_  = \new_Sorter100|6568_  & \new_Sorter100|6569_ ;
  assign \new_Sorter100|6669_  = \new_Sorter100|6568_  | \new_Sorter100|6569_ ;
  assign \new_Sorter100|6670_  = \new_Sorter100|6570_  & \new_Sorter100|6571_ ;
  assign \new_Sorter100|6671_  = \new_Sorter100|6570_  | \new_Sorter100|6571_ ;
  assign \new_Sorter100|6672_  = \new_Sorter100|6572_  & \new_Sorter100|6573_ ;
  assign \new_Sorter100|6673_  = \new_Sorter100|6572_  | \new_Sorter100|6573_ ;
  assign \new_Sorter100|6674_  = \new_Sorter100|6574_  & \new_Sorter100|6575_ ;
  assign \new_Sorter100|6675_  = \new_Sorter100|6574_  | \new_Sorter100|6575_ ;
  assign \new_Sorter100|6676_  = \new_Sorter100|6576_  & \new_Sorter100|6577_ ;
  assign \new_Sorter100|6677_  = \new_Sorter100|6576_  | \new_Sorter100|6577_ ;
  assign \new_Sorter100|6678_  = \new_Sorter100|6578_  & \new_Sorter100|6579_ ;
  assign \new_Sorter100|6679_  = \new_Sorter100|6578_  | \new_Sorter100|6579_ ;
  assign \new_Sorter100|6680_  = \new_Sorter100|6580_  & \new_Sorter100|6581_ ;
  assign \new_Sorter100|6681_  = \new_Sorter100|6580_  | \new_Sorter100|6581_ ;
  assign \new_Sorter100|6682_  = \new_Sorter100|6582_  & \new_Sorter100|6583_ ;
  assign \new_Sorter100|6683_  = \new_Sorter100|6582_  | \new_Sorter100|6583_ ;
  assign \new_Sorter100|6684_  = \new_Sorter100|6584_  & \new_Sorter100|6585_ ;
  assign \new_Sorter100|6685_  = \new_Sorter100|6584_  | \new_Sorter100|6585_ ;
  assign \new_Sorter100|6686_  = \new_Sorter100|6586_  & \new_Sorter100|6587_ ;
  assign \new_Sorter100|6687_  = \new_Sorter100|6586_  | \new_Sorter100|6587_ ;
  assign \new_Sorter100|6688_  = \new_Sorter100|6588_  & \new_Sorter100|6589_ ;
  assign \new_Sorter100|6689_  = \new_Sorter100|6588_  | \new_Sorter100|6589_ ;
  assign \new_Sorter100|6690_  = \new_Sorter100|6590_  & \new_Sorter100|6591_ ;
  assign \new_Sorter100|6691_  = \new_Sorter100|6590_  | \new_Sorter100|6591_ ;
  assign \new_Sorter100|6692_  = \new_Sorter100|6592_  & \new_Sorter100|6593_ ;
  assign \new_Sorter100|6693_  = \new_Sorter100|6592_  | \new_Sorter100|6593_ ;
  assign \new_Sorter100|6694_  = \new_Sorter100|6594_  & \new_Sorter100|6595_ ;
  assign \new_Sorter100|6695_  = \new_Sorter100|6594_  | \new_Sorter100|6595_ ;
  assign \new_Sorter100|6696_  = \new_Sorter100|6596_  & \new_Sorter100|6597_ ;
  assign \new_Sorter100|6697_  = \new_Sorter100|6596_  | \new_Sorter100|6597_ ;
  assign \new_Sorter100|6698_  = \new_Sorter100|6598_  & \new_Sorter100|6599_ ;
  assign \new_Sorter100|6699_  = \new_Sorter100|6598_  | \new_Sorter100|6599_ ;
  assign \new_Sorter100|6700_  = \new_Sorter100|6600_ ;
  assign \new_Sorter100|6799_  = \new_Sorter100|6699_ ;
  assign \new_Sorter100|6701_  = \new_Sorter100|6601_  & \new_Sorter100|6602_ ;
  assign \new_Sorter100|6702_  = \new_Sorter100|6601_  | \new_Sorter100|6602_ ;
  assign \new_Sorter100|6703_  = \new_Sorter100|6603_  & \new_Sorter100|6604_ ;
  assign \new_Sorter100|6704_  = \new_Sorter100|6603_  | \new_Sorter100|6604_ ;
  assign \new_Sorter100|6705_  = \new_Sorter100|6605_  & \new_Sorter100|6606_ ;
  assign \new_Sorter100|6706_  = \new_Sorter100|6605_  | \new_Sorter100|6606_ ;
  assign \new_Sorter100|6707_  = \new_Sorter100|6607_  & \new_Sorter100|6608_ ;
  assign \new_Sorter100|6708_  = \new_Sorter100|6607_  | \new_Sorter100|6608_ ;
  assign \new_Sorter100|6709_  = \new_Sorter100|6609_  & \new_Sorter100|6610_ ;
  assign \new_Sorter100|6710_  = \new_Sorter100|6609_  | \new_Sorter100|6610_ ;
  assign \new_Sorter100|6711_  = \new_Sorter100|6611_  & \new_Sorter100|6612_ ;
  assign \new_Sorter100|6712_  = \new_Sorter100|6611_  | \new_Sorter100|6612_ ;
  assign \new_Sorter100|6713_  = \new_Sorter100|6613_  & \new_Sorter100|6614_ ;
  assign \new_Sorter100|6714_  = \new_Sorter100|6613_  | \new_Sorter100|6614_ ;
  assign \new_Sorter100|6715_  = \new_Sorter100|6615_  & \new_Sorter100|6616_ ;
  assign \new_Sorter100|6716_  = \new_Sorter100|6615_  | \new_Sorter100|6616_ ;
  assign \new_Sorter100|6717_  = \new_Sorter100|6617_  & \new_Sorter100|6618_ ;
  assign \new_Sorter100|6718_  = \new_Sorter100|6617_  | \new_Sorter100|6618_ ;
  assign \new_Sorter100|6719_  = \new_Sorter100|6619_  & \new_Sorter100|6620_ ;
  assign \new_Sorter100|6720_  = \new_Sorter100|6619_  | \new_Sorter100|6620_ ;
  assign \new_Sorter100|6721_  = \new_Sorter100|6621_  & \new_Sorter100|6622_ ;
  assign \new_Sorter100|6722_  = \new_Sorter100|6621_  | \new_Sorter100|6622_ ;
  assign \new_Sorter100|6723_  = \new_Sorter100|6623_  & \new_Sorter100|6624_ ;
  assign \new_Sorter100|6724_  = \new_Sorter100|6623_  | \new_Sorter100|6624_ ;
  assign \new_Sorter100|6725_  = \new_Sorter100|6625_  & \new_Sorter100|6626_ ;
  assign \new_Sorter100|6726_  = \new_Sorter100|6625_  | \new_Sorter100|6626_ ;
  assign \new_Sorter100|6727_  = \new_Sorter100|6627_  & \new_Sorter100|6628_ ;
  assign \new_Sorter100|6728_  = \new_Sorter100|6627_  | \new_Sorter100|6628_ ;
  assign \new_Sorter100|6729_  = \new_Sorter100|6629_  & \new_Sorter100|6630_ ;
  assign \new_Sorter100|6730_  = \new_Sorter100|6629_  | \new_Sorter100|6630_ ;
  assign \new_Sorter100|6731_  = \new_Sorter100|6631_  & \new_Sorter100|6632_ ;
  assign \new_Sorter100|6732_  = \new_Sorter100|6631_  | \new_Sorter100|6632_ ;
  assign \new_Sorter100|6733_  = \new_Sorter100|6633_  & \new_Sorter100|6634_ ;
  assign \new_Sorter100|6734_  = \new_Sorter100|6633_  | \new_Sorter100|6634_ ;
  assign \new_Sorter100|6735_  = \new_Sorter100|6635_  & \new_Sorter100|6636_ ;
  assign \new_Sorter100|6736_  = \new_Sorter100|6635_  | \new_Sorter100|6636_ ;
  assign \new_Sorter100|6737_  = \new_Sorter100|6637_  & \new_Sorter100|6638_ ;
  assign \new_Sorter100|6738_  = \new_Sorter100|6637_  | \new_Sorter100|6638_ ;
  assign \new_Sorter100|6739_  = \new_Sorter100|6639_  & \new_Sorter100|6640_ ;
  assign \new_Sorter100|6740_  = \new_Sorter100|6639_  | \new_Sorter100|6640_ ;
  assign \new_Sorter100|6741_  = \new_Sorter100|6641_  & \new_Sorter100|6642_ ;
  assign \new_Sorter100|6742_  = \new_Sorter100|6641_  | \new_Sorter100|6642_ ;
  assign \new_Sorter100|6743_  = \new_Sorter100|6643_  & \new_Sorter100|6644_ ;
  assign \new_Sorter100|6744_  = \new_Sorter100|6643_  | \new_Sorter100|6644_ ;
  assign \new_Sorter100|6745_  = \new_Sorter100|6645_  & \new_Sorter100|6646_ ;
  assign \new_Sorter100|6746_  = \new_Sorter100|6645_  | \new_Sorter100|6646_ ;
  assign \new_Sorter100|6747_  = \new_Sorter100|6647_  & \new_Sorter100|6648_ ;
  assign \new_Sorter100|6748_  = \new_Sorter100|6647_  | \new_Sorter100|6648_ ;
  assign \new_Sorter100|6749_  = \new_Sorter100|6649_  & \new_Sorter100|6650_ ;
  assign \new_Sorter100|6750_  = \new_Sorter100|6649_  | \new_Sorter100|6650_ ;
  assign \new_Sorter100|6751_  = \new_Sorter100|6651_  & \new_Sorter100|6652_ ;
  assign \new_Sorter100|6752_  = \new_Sorter100|6651_  | \new_Sorter100|6652_ ;
  assign \new_Sorter100|6753_  = \new_Sorter100|6653_  & \new_Sorter100|6654_ ;
  assign \new_Sorter100|6754_  = \new_Sorter100|6653_  | \new_Sorter100|6654_ ;
  assign \new_Sorter100|6755_  = \new_Sorter100|6655_  & \new_Sorter100|6656_ ;
  assign \new_Sorter100|6756_  = \new_Sorter100|6655_  | \new_Sorter100|6656_ ;
  assign \new_Sorter100|6757_  = \new_Sorter100|6657_  & \new_Sorter100|6658_ ;
  assign \new_Sorter100|6758_  = \new_Sorter100|6657_  | \new_Sorter100|6658_ ;
  assign \new_Sorter100|6759_  = \new_Sorter100|6659_  & \new_Sorter100|6660_ ;
  assign \new_Sorter100|6760_  = \new_Sorter100|6659_  | \new_Sorter100|6660_ ;
  assign \new_Sorter100|6761_  = \new_Sorter100|6661_  & \new_Sorter100|6662_ ;
  assign \new_Sorter100|6762_  = \new_Sorter100|6661_  | \new_Sorter100|6662_ ;
  assign \new_Sorter100|6763_  = \new_Sorter100|6663_  & \new_Sorter100|6664_ ;
  assign \new_Sorter100|6764_  = \new_Sorter100|6663_  | \new_Sorter100|6664_ ;
  assign \new_Sorter100|6765_  = \new_Sorter100|6665_  & \new_Sorter100|6666_ ;
  assign \new_Sorter100|6766_  = \new_Sorter100|6665_  | \new_Sorter100|6666_ ;
  assign \new_Sorter100|6767_  = \new_Sorter100|6667_  & \new_Sorter100|6668_ ;
  assign \new_Sorter100|6768_  = \new_Sorter100|6667_  | \new_Sorter100|6668_ ;
  assign \new_Sorter100|6769_  = \new_Sorter100|6669_  & \new_Sorter100|6670_ ;
  assign \new_Sorter100|6770_  = \new_Sorter100|6669_  | \new_Sorter100|6670_ ;
  assign \new_Sorter100|6771_  = \new_Sorter100|6671_  & \new_Sorter100|6672_ ;
  assign \new_Sorter100|6772_  = \new_Sorter100|6671_  | \new_Sorter100|6672_ ;
  assign \new_Sorter100|6773_  = \new_Sorter100|6673_  & \new_Sorter100|6674_ ;
  assign \new_Sorter100|6774_  = \new_Sorter100|6673_  | \new_Sorter100|6674_ ;
  assign \new_Sorter100|6775_  = \new_Sorter100|6675_  & \new_Sorter100|6676_ ;
  assign \new_Sorter100|6776_  = \new_Sorter100|6675_  | \new_Sorter100|6676_ ;
  assign \new_Sorter100|6777_  = \new_Sorter100|6677_  & \new_Sorter100|6678_ ;
  assign \new_Sorter100|6778_  = \new_Sorter100|6677_  | \new_Sorter100|6678_ ;
  assign \new_Sorter100|6779_  = \new_Sorter100|6679_  & \new_Sorter100|6680_ ;
  assign \new_Sorter100|6780_  = \new_Sorter100|6679_  | \new_Sorter100|6680_ ;
  assign \new_Sorter100|6781_  = \new_Sorter100|6681_  & \new_Sorter100|6682_ ;
  assign \new_Sorter100|6782_  = \new_Sorter100|6681_  | \new_Sorter100|6682_ ;
  assign \new_Sorter100|6783_  = \new_Sorter100|6683_  & \new_Sorter100|6684_ ;
  assign \new_Sorter100|6784_  = \new_Sorter100|6683_  | \new_Sorter100|6684_ ;
  assign \new_Sorter100|6785_  = \new_Sorter100|6685_  & \new_Sorter100|6686_ ;
  assign \new_Sorter100|6786_  = \new_Sorter100|6685_  | \new_Sorter100|6686_ ;
  assign \new_Sorter100|6787_  = \new_Sorter100|6687_  & \new_Sorter100|6688_ ;
  assign \new_Sorter100|6788_  = \new_Sorter100|6687_  | \new_Sorter100|6688_ ;
  assign \new_Sorter100|6789_  = \new_Sorter100|6689_  & \new_Sorter100|6690_ ;
  assign \new_Sorter100|6790_  = \new_Sorter100|6689_  | \new_Sorter100|6690_ ;
  assign \new_Sorter100|6791_  = \new_Sorter100|6691_  & \new_Sorter100|6692_ ;
  assign \new_Sorter100|6792_  = \new_Sorter100|6691_  | \new_Sorter100|6692_ ;
  assign \new_Sorter100|6793_  = \new_Sorter100|6693_  & \new_Sorter100|6694_ ;
  assign \new_Sorter100|6794_  = \new_Sorter100|6693_  | \new_Sorter100|6694_ ;
  assign \new_Sorter100|6795_  = \new_Sorter100|6695_  & \new_Sorter100|6696_ ;
  assign \new_Sorter100|6796_  = \new_Sorter100|6695_  | \new_Sorter100|6696_ ;
  assign \new_Sorter100|6797_  = \new_Sorter100|6697_  & \new_Sorter100|6698_ ;
  assign \new_Sorter100|6798_  = \new_Sorter100|6697_  | \new_Sorter100|6698_ ;
  assign \new_Sorter100|6800_  = \new_Sorter100|6700_  & \new_Sorter100|6701_ ;
  assign \new_Sorter100|6801_  = \new_Sorter100|6700_  | \new_Sorter100|6701_ ;
  assign \new_Sorter100|6802_  = \new_Sorter100|6702_  & \new_Sorter100|6703_ ;
  assign \new_Sorter100|6803_  = \new_Sorter100|6702_  | \new_Sorter100|6703_ ;
  assign \new_Sorter100|6804_  = \new_Sorter100|6704_  & \new_Sorter100|6705_ ;
  assign \new_Sorter100|6805_  = \new_Sorter100|6704_  | \new_Sorter100|6705_ ;
  assign \new_Sorter100|6806_  = \new_Sorter100|6706_  & \new_Sorter100|6707_ ;
  assign \new_Sorter100|6807_  = \new_Sorter100|6706_  | \new_Sorter100|6707_ ;
  assign \new_Sorter100|6808_  = \new_Sorter100|6708_  & \new_Sorter100|6709_ ;
  assign \new_Sorter100|6809_  = \new_Sorter100|6708_  | \new_Sorter100|6709_ ;
  assign \new_Sorter100|6810_  = \new_Sorter100|6710_  & \new_Sorter100|6711_ ;
  assign \new_Sorter100|6811_  = \new_Sorter100|6710_  | \new_Sorter100|6711_ ;
  assign \new_Sorter100|6812_  = \new_Sorter100|6712_  & \new_Sorter100|6713_ ;
  assign \new_Sorter100|6813_  = \new_Sorter100|6712_  | \new_Sorter100|6713_ ;
  assign \new_Sorter100|6814_  = \new_Sorter100|6714_  & \new_Sorter100|6715_ ;
  assign \new_Sorter100|6815_  = \new_Sorter100|6714_  | \new_Sorter100|6715_ ;
  assign \new_Sorter100|6816_  = \new_Sorter100|6716_  & \new_Sorter100|6717_ ;
  assign \new_Sorter100|6817_  = \new_Sorter100|6716_  | \new_Sorter100|6717_ ;
  assign \new_Sorter100|6818_  = \new_Sorter100|6718_  & \new_Sorter100|6719_ ;
  assign \new_Sorter100|6819_  = \new_Sorter100|6718_  | \new_Sorter100|6719_ ;
  assign \new_Sorter100|6820_  = \new_Sorter100|6720_  & \new_Sorter100|6721_ ;
  assign \new_Sorter100|6821_  = \new_Sorter100|6720_  | \new_Sorter100|6721_ ;
  assign \new_Sorter100|6822_  = \new_Sorter100|6722_  & \new_Sorter100|6723_ ;
  assign \new_Sorter100|6823_  = \new_Sorter100|6722_  | \new_Sorter100|6723_ ;
  assign \new_Sorter100|6824_  = \new_Sorter100|6724_  & \new_Sorter100|6725_ ;
  assign \new_Sorter100|6825_  = \new_Sorter100|6724_  | \new_Sorter100|6725_ ;
  assign \new_Sorter100|6826_  = \new_Sorter100|6726_  & \new_Sorter100|6727_ ;
  assign \new_Sorter100|6827_  = \new_Sorter100|6726_  | \new_Sorter100|6727_ ;
  assign \new_Sorter100|6828_  = \new_Sorter100|6728_  & \new_Sorter100|6729_ ;
  assign \new_Sorter100|6829_  = \new_Sorter100|6728_  | \new_Sorter100|6729_ ;
  assign \new_Sorter100|6830_  = \new_Sorter100|6730_  & \new_Sorter100|6731_ ;
  assign \new_Sorter100|6831_  = \new_Sorter100|6730_  | \new_Sorter100|6731_ ;
  assign \new_Sorter100|6832_  = \new_Sorter100|6732_  & \new_Sorter100|6733_ ;
  assign \new_Sorter100|6833_  = \new_Sorter100|6732_  | \new_Sorter100|6733_ ;
  assign \new_Sorter100|6834_  = \new_Sorter100|6734_  & \new_Sorter100|6735_ ;
  assign \new_Sorter100|6835_  = \new_Sorter100|6734_  | \new_Sorter100|6735_ ;
  assign \new_Sorter100|6836_  = \new_Sorter100|6736_  & \new_Sorter100|6737_ ;
  assign \new_Sorter100|6837_  = \new_Sorter100|6736_  | \new_Sorter100|6737_ ;
  assign \new_Sorter100|6838_  = \new_Sorter100|6738_  & \new_Sorter100|6739_ ;
  assign \new_Sorter100|6839_  = \new_Sorter100|6738_  | \new_Sorter100|6739_ ;
  assign \new_Sorter100|6840_  = \new_Sorter100|6740_  & \new_Sorter100|6741_ ;
  assign \new_Sorter100|6841_  = \new_Sorter100|6740_  | \new_Sorter100|6741_ ;
  assign \new_Sorter100|6842_  = \new_Sorter100|6742_  & \new_Sorter100|6743_ ;
  assign \new_Sorter100|6843_  = \new_Sorter100|6742_  | \new_Sorter100|6743_ ;
  assign \new_Sorter100|6844_  = \new_Sorter100|6744_  & \new_Sorter100|6745_ ;
  assign \new_Sorter100|6845_  = \new_Sorter100|6744_  | \new_Sorter100|6745_ ;
  assign \new_Sorter100|6846_  = \new_Sorter100|6746_  & \new_Sorter100|6747_ ;
  assign \new_Sorter100|6847_  = \new_Sorter100|6746_  | \new_Sorter100|6747_ ;
  assign \new_Sorter100|6848_  = \new_Sorter100|6748_  & \new_Sorter100|6749_ ;
  assign \new_Sorter100|6849_  = \new_Sorter100|6748_  | \new_Sorter100|6749_ ;
  assign \new_Sorter100|6850_  = \new_Sorter100|6750_  & \new_Sorter100|6751_ ;
  assign \new_Sorter100|6851_  = \new_Sorter100|6750_  | \new_Sorter100|6751_ ;
  assign \new_Sorter100|6852_  = \new_Sorter100|6752_  & \new_Sorter100|6753_ ;
  assign \new_Sorter100|6853_  = \new_Sorter100|6752_  | \new_Sorter100|6753_ ;
  assign \new_Sorter100|6854_  = \new_Sorter100|6754_  & \new_Sorter100|6755_ ;
  assign \new_Sorter100|6855_  = \new_Sorter100|6754_  | \new_Sorter100|6755_ ;
  assign \new_Sorter100|6856_  = \new_Sorter100|6756_  & \new_Sorter100|6757_ ;
  assign \new_Sorter100|6857_  = \new_Sorter100|6756_  | \new_Sorter100|6757_ ;
  assign \new_Sorter100|6858_  = \new_Sorter100|6758_  & \new_Sorter100|6759_ ;
  assign \new_Sorter100|6859_  = \new_Sorter100|6758_  | \new_Sorter100|6759_ ;
  assign \new_Sorter100|6860_  = \new_Sorter100|6760_  & \new_Sorter100|6761_ ;
  assign \new_Sorter100|6861_  = \new_Sorter100|6760_  | \new_Sorter100|6761_ ;
  assign \new_Sorter100|6862_  = \new_Sorter100|6762_  & \new_Sorter100|6763_ ;
  assign \new_Sorter100|6863_  = \new_Sorter100|6762_  | \new_Sorter100|6763_ ;
  assign \new_Sorter100|6864_  = \new_Sorter100|6764_  & \new_Sorter100|6765_ ;
  assign \new_Sorter100|6865_  = \new_Sorter100|6764_  | \new_Sorter100|6765_ ;
  assign \new_Sorter100|6866_  = \new_Sorter100|6766_  & \new_Sorter100|6767_ ;
  assign \new_Sorter100|6867_  = \new_Sorter100|6766_  | \new_Sorter100|6767_ ;
  assign \new_Sorter100|6868_  = \new_Sorter100|6768_  & \new_Sorter100|6769_ ;
  assign \new_Sorter100|6869_  = \new_Sorter100|6768_  | \new_Sorter100|6769_ ;
  assign \new_Sorter100|6870_  = \new_Sorter100|6770_  & \new_Sorter100|6771_ ;
  assign \new_Sorter100|6871_  = \new_Sorter100|6770_  | \new_Sorter100|6771_ ;
  assign \new_Sorter100|6872_  = \new_Sorter100|6772_  & \new_Sorter100|6773_ ;
  assign \new_Sorter100|6873_  = \new_Sorter100|6772_  | \new_Sorter100|6773_ ;
  assign \new_Sorter100|6874_  = \new_Sorter100|6774_  & \new_Sorter100|6775_ ;
  assign \new_Sorter100|6875_  = \new_Sorter100|6774_  | \new_Sorter100|6775_ ;
  assign \new_Sorter100|6876_  = \new_Sorter100|6776_  & \new_Sorter100|6777_ ;
  assign \new_Sorter100|6877_  = \new_Sorter100|6776_  | \new_Sorter100|6777_ ;
  assign \new_Sorter100|6878_  = \new_Sorter100|6778_  & \new_Sorter100|6779_ ;
  assign \new_Sorter100|6879_  = \new_Sorter100|6778_  | \new_Sorter100|6779_ ;
  assign \new_Sorter100|6880_  = \new_Sorter100|6780_  & \new_Sorter100|6781_ ;
  assign \new_Sorter100|6881_  = \new_Sorter100|6780_  | \new_Sorter100|6781_ ;
  assign \new_Sorter100|6882_  = \new_Sorter100|6782_  & \new_Sorter100|6783_ ;
  assign \new_Sorter100|6883_  = \new_Sorter100|6782_  | \new_Sorter100|6783_ ;
  assign \new_Sorter100|6884_  = \new_Sorter100|6784_  & \new_Sorter100|6785_ ;
  assign \new_Sorter100|6885_  = \new_Sorter100|6784_  | \new_Sorter100|6785_ ;
  assign \new_Sorter100|6886_  = \new_Sorter100|6786_  & \new_Sorter100|6787_ ;
  assign \new_Sorter100|6887_  = \new_Sorter100|6786_  | \new_Sorter100|6787_ ;
  assign \new_Sorter100|6888_  = \new_Sorter100|6788_  & \new_Sorter100|6789_ ;
  assign \new_Sorter100|6889_  = \new_Sorter100|6788_  | \new_Sorter100|6789_ ;
  assign \new_Sorter100|6890_  = \new_Sorter100|6790_  & \new_Sorter100|6791_ ;
  assign \new_Sorter100|6891_  = \new_Sorter100|6790_  | \new_Sorter100|6791_ ;
  assign \new_Sorter100|6892_  = \new_Sorter100|6792_  & \new_Sorter100|6793_ ;
  assign \new_Sorter100|6893_  = \new_Sorter100|6792_  | \new_Sorter100|6793_ ;
  assign \new_Sorter100|6894_  = \new_Sorter100|6794_  & \new_Sorter100|6795_ ;
  assign \new_Sorter100|6895_  = \new_Sorter100|6794_  | \new_Sorter100|6795_ ;
  assign \new_Sorter100|6896_  = \new_Sorter100|6796_  & \new_Sorter100|6797_ ;
  assign \new_Sorter100|6897_  = \new_Sorter100|6796_  | \new_Sorter100|6797_ ;
  assign \new_Sorter100|6898_  = \new_Sorter100|6798_  & \new_Sorter100|6799_ ;
  assign \new_Sorter100|6899_  = \new_Sorter100|6798_  | \new_Sorter100|6799_ ;
  assign \new_Sorter100|6900_  = \new_Sorter100|6800_ ;
  assign \new_Sorter100|6999_  = \new_Sorter100|6899_ ;
  assign \new_Sorter100|6901_  = \new_Sorter100|6801_  & \new_Sorter100|6802_ ;
  assign \new_Sorter100|6902_  = \new_Sorter100|6801_  | \new_Sorter100|6802_ ;
  assign \new_Sorter100|6903_  = \new_Sorter100|6803_  & \new_Sorter100|6804_ ;
  assign \new_Sorter100|6904_  = \new_Sorter100|6803_  | \new_Sorter100|6804_ ;
  assign \new_Sorter100|6905_  = \new_Sorter100|6805_  & \new_Sorter100|6806_ ;
  assign \new_Sorter100|6906_  = \new_Sorter100|6805_  | \new_Sorter100|6806_ ;
  assign \new_Sorter100|6907_  = \new_Sorter100|6807_  & \new_Sorter100|6808_ ;
  assign \new_Sorter100|6908_  = \new_Sorter100|6807_  | \new_Sorter100|6808_ ;
  assign \new_Sorter100|6909_  = \new_Sorter100|6809_  & \new_Sorter100|6810_ ;
  assign \new_Sorter100|6910_  = \new_Sorter100|6809_  | \new_Sorter100|6810_ ;
  assign \new_Sorter100|6911_  = \new_Sorter100|6811_  & \new_Sorter100|6812_ ;
  assign \new_Sorter100|6912_  = \new_Sorter100|6811_  | \new_Sorter100|6812_ ;
  assign \new_Sorter100|6913_  = \new_Sorter100|6813_  & \new_Sorter100|6814_ ;
  assign \new_Sorter100|6914_  = \new_Sorter100|6813_  | \new_Sorter100|6814_ ;
  assign \new_Sorter100|6915_  = \new_Sorter100|6815_  & \new_Sorter100|6816_ ;
  assign \new_Sorter100|6916_  = \new_Sorter100|6815_  | \new_Sorter100|6816_ ;
  assign \new_Sorter100|6917_  = \new_Sorter100|6817_  & \new_Sorter100|6818_ ;
  assign \new_Sorter100|6918_  = \new_Sorter100|6817_  | \new_Sorter100|6818_ ;
  assign \new_Sorter100|6919_  = \new_Sorter100|6819_  & \new_Sorter100|6820_ ;
  assign \new_Sorter100|6920_  = \new_Sorter100|6819_  | \new_Sorter100|6820_ ;
  assign \new_Sorter100|6921_  = \new_Sorter100|6821_  & \new_Sorter100|6822_ ;
  assign \new_Sorter100|6922_  = \new_Sorter100|6821_  | \new_Sorter100|6822_ ;
  assign \new_Sorter100|6923_  = \new_Sorter100|6823_  & \new_Sorter100|6824_ ;
  assign \new_Sorter100|6924_  = \new_Sorter100|6823_  | \new_Sorter100|6824_ ;
  assign \new_Sorter100|6925_  = \new_Sorter100|6825_  & \new_Sorter100|6826_ ;
  assign \new_Sorter100|6926_  = \new_Sorter100|6825_  | \new_Sorter100|6826_ ;
  assign \new_Sorter100|6927_  = \new_Sorter100|6827_  & \new_Sorter100|6828_ ;
  assign \new_Sorter100|6928_  = \new_Sorter100|6827_  | \new_Sorter100|6828_ ;
  assign \new_Sorter100|6929_  = \new_Sorter100|6829_  & \new_Sorter100|6830_ ;
  assign \new_Sorter100|6930_  = \new_Sorter100|6829_  | \new_Sorter100|6830_ ;
  assign \new_Sorter100|6931_  = \new_Sorter100|6831_  & \new_Sorter100|6832_ ;
  assign \new_Sorter100|6932_  = \new_Sorter100|6831_  | \new_Sorter100|6832_ ;
  assign \new_Sorter100|6933_  = \new_Sorter100|6833_  & \new_Sorter100|6834_ ;
  assign \new_Sorter100|6934_  = \new_Sorter100|6833_  | \new_Sorter100|6834_ ;
  assign \new_Sorter100|6935_  = \new_Sorter100|6835_  & \new_Sorter100|6836_ ;
  assign \new_Sorter100|6936_  = \new_Sorter100|6835_  | \new_Sorter100|6836_ ;
  assign \new_Sorter100|6937_  = \new_Sorter100|6837_  & \new_Sorter100|6838_ ;
  assign \new_Sorter100|6938_  = \new_Sorter100|6837_  | \new_Sorter100|6838_ ;
  assign \new_Sorter100|6939_  = \new_Sorter100|6839_  & \new_Sorter100|6840_ ;
  assign \new_Sorter100|6940_  = \new_Sorter100|6839_  | \new_Sorter100|6840_ ;
  assign \new_Sorter100|6941_  = \new_Sorter100|6841_  & \new_Sorter100|6842_ ;
  assign \new_Sorter100|6942_  = \new_Sorter100|6841_  | \new_Sorter100|6842_ ;
  assign \new_Sorter100|6943_  = \new_Sorter100|6843_  & \new_Sorter100|6844_ ;
  assign \new_Sorter100|6944_  = \new_Sorter100|6843_  | \new_Sorter100|6844_ ;
  assign \new_Sorter100|6945_  = \new_Sorter100|6845_  & \new_Sorter100|6846_ ;
  assign \new_Sorter100|6946_  = \new_Sorter100|6845_  | \new_Sorter100|6846_ ;
  assign \new_Sorter100|6947_  = \new_Sorter100|6847_  & \new_Sorter100|6848_ ;
  assign \new_Sorter100|6948_  = \new_Sorter100|6847_  | \new_Sorter100|6848_ ;
  assign \new_Sorter100|6949_  = \new_Sorter100|6849_  & \new_Sorter100|6850_ ;
  assign \new_Sorter100|6950_  = \new_Sorter100|6849_  | \new_Sorter100|6850_ ;
  assign \new_Sorter100|6951_  = \new_Sorter100|6851_  & \new_Sorter100|6852_ ;
  assign \new_Sorter100|6952_  = \new_Sorter100|6851_  | \new_Sorter100|6852_ ;
  assign \new_Sorter100|6953_  = \new_Sorter100|6853_  & \new_Sorter100|6854_ ;
  assign \new_Sorter100|6954_  = \new_Sorter100|6853_  | \new_Sorter100|6854_ ;
  assign \new_Sorter100|6955_  = \new_Sorter100|6855_  & \new_Sorter100|6856_ ;
  assign \new_Sorter100|6956_  = \new_Sorter100|6855_  | \new_Sorter100|6856_ ;
  assign \new_Sorter100|6957_  = \new_Sorter100|6857_  & \new_Sorter100|6858_ ;
  assign \new_Sorter100|6958_  = \new_Sorter100|6857_  | \new_Sorter100|6858_ ;
  assign \new_Sorter100|6959_  = \new_Sorter100|6859_  & \new_Sorter100|6860_ ;
  assign \new_Sorter100|6960_  = \new_Sorter100|6859_  | \new_Sorter100|6860_ ;
  assign \new_Sorter100|6961_  = \new_Sorter100|6861_  & \new_Sorter100|6862_ ;
  assign \new_Sorter100|6962_  = \new_Sorter100|6861_  | \new_Sorter100|6862_ ;
  assign \new_Sorter100|6963_  = \new_Sorter100|6863_  & \new_Sorter100|6864_ ;
  assign \new_Sorter100|6964_  = \new_Sorter100|6863_  | \new_Sorter100|6864_ ;
  assign \new_Sorter100|6965_  = \new_Sorter100|6865_  & \new_Sorter100|6866_ ;
  assign \new_Sorter100|6966_  = \new_Sorter100|6865_  | \new_Sorter100|6866_ ;
  assign \new_Sorter100|6967_  = \new_Sorter100|6867_  & \new_Sorter100|6868_ ;
  assign \new_Sorter100|6968_  = \new_Sorter100|6867_  | \new_Sorter100|6868_ ;
  assign \new_Sorter100|6969_  = \new_Sorter100|6869_  & \new_Sorter100|6870_ ;
  assign \new_Sorter100|6970_  = \new_Sorter100|6869_  | \new_Sorter100|6870_ ;
  assign \new_Sorter100|6971_  = \new_Sorter100|6871_  & \new_Sorter100|6872_ ;
  assign \new_Sorter100|6972_  = \new_Sorter100|6871_  | \new_Sorter100|6872_ ;
  assign \new_Sorter100|6973_  = \new_Sorter100|6873_  & \new_Sorter100|6874_ ;
  assign \new_Sorter100|6974_  = \new_Sorter100|6873_  | \new_Sorter100|6874_ ;
  assign \new_Sorter100|6975_  = \new_Sorter100|6875_  & \new_Sorter100|6876_ ;
  assign \new_Sorter100|6976_  = \new_Sorter100|6875_  | \new_Sorter100|6876_ ;
  assign \new_Sorter100|6977_  = \new_Sorter100|6877_  & \new_Sorter100|6878_ ;
  assign \new_Sorter100|6978_  = \new_Sorter100|6877_  | \new_Sorter100|6878_ ;
  assign \new_Sorter100|6979_  = \new_Sorter100|6879_  & \new_Sorter100|6880_ ;
  assign \new_Sorter100|6980_  = \new_Sorter100|6879_  | \new_Sorter100|6880_ ;
  assign \new_Sorter100|6981_  = \new_Sorter100|6881_  & \new_Sorter100|6882_ ;
  assign \new_Sorter100|6982_  = \new_Sorter100|6881_  | \new_Sorter100|6882_ ;
  assign \new_Sorter100|6983_  = \new_Sorter100|6883_  & \new_Sorter100|6884_ ;
  assign \new_Sorter100|6984_  = \new_Sorter100|6883_  | \new_Sorter100|6884_ ;
  assign \new_Sorter100|6985_  = \new_Sorter100|6885_  & \new_Sorter100|6886_ ;
  assign \new_Sorter100|6986_  = \new_Sorter100|6885_  | \new_Sorter100|6886_ ;
  assign \new_Sorter100|6987_  = \new_Sorter100|6887_  & \new_Sorter100|6888_ ;
  assign \new_Sorter100|6988_  = \new_Sorter100|6887_  | \new_Sorter100|6888_ ;
  assign \new_Sorter100|6989_  = \new_Sorter100|6889_  & \new_Sorter100|6890_ ;
  assign \new_Sorter100|6990_  = \new_Sorter100|6889_  | \new_Sorter100|6890_ ;
  assign \new_Sorter100|6991_  = \new_Sorter100|6891_  & \new_Sorter100|6892_ ;
  assign \new_Sorter100|6992_  = \new_Sorter100|6891_  | \new_Sorter100|6892_ ;
  assign \new_Sorter100|6993_  = \new_Sorter100|6893_  & \new_Sorter100|6894_ ;
  assign \new_Sorter100|6994_  = \new_Sorter100|6893_  | \new_Sorter100|6894_ ;
  assign \new_Sorter100|6995_  = \new_Sorter100|6895_  & \new_Sorter100|6896_ ;
  assign \new_Sorter100|6996_  = \new_Sorter100|6895_  | \new_Sorter100|6896_ ;
  assign \new_Sorter100|6997_  = \new_Sorter100|6897_  & \new_Sorter100|6898_ ;
  assign \new_Sorter100|6998_  = \new_Sorter100|6897_  | \new_Sorter100|6898_ ;
  assign \new_Sorter100|7000_  = \new_Sorter100|6900_  & \new_Sorter100|6901_ ;
  assign \new_Sorter100|7001_  = \new_Sorter100|6900_  | \new_Sorter100|6901_ ;
  assign \new_Sorter100|7002_  = \new_Sorter100|6902_  & \new_Sorter100|6903_ ;
  assign \new_Sorter100|7003_  = \new_Sorter100|6902_  | \new_Sorter100|6903_ ;
  assign \new_Sorter100|7004_  = \new_Sorter100|6904_  & \new_Sorter100|6905_ ;
  assign \new_Sorter100|7005_  = \new_Sorter100|6904_  | \new_Sorter100|6905_ ;
  assign \new_Sorter100|7006_  = \new_Sorter100|6906_  & \new_Sorter100|6907_ ;
  assign \new_Sorter100|7007_  = \new_Sorter100|6906_  | \new_Sorter100|6907_ ;
  assign \new_Sorter100|7008_  = \new_Sorter100|6908_  & \new_Sorter100|6909_ ;
  assign \new_Sorter100|7009_  = \new_Sorter100|6908_  | \new_Sorter100|6909_ ;
  assign \new_Sorter100|7010_  = \new_Sorter100|6910_  & \new_Sorter100|6911_ ;
  assign \new_Sorter100|7011_  = \new_Sorter100|6910_  | \new_Sorter100|6911_ ;
  assign \new_Sorter100|7012_  = \new_Sorter100|6912_  & \new_Sorter100|6913_ ;
  assign \new_Sorter100|7013_  = \new_Sorter100|6912_  | \new_Sorter100|6913_ ;
  assign \new_Sorter100|7014_  = \new_Sorter100|6914_  & \new_Sorter100|6915_ ;
  assign \new_Sorter100|7015_  = \new_Sorter100|6914_  | \new_Sorter100|6915_ ;
  assign \new_Sorter100|7016_  = \new_Sorter100|6916_  & \new_Sorter100|6917_ ;
  assign \new_Sorter100|7017_  = \new_Sorter100|6916_  | \new_Sorter100|6917_ ;
  assign \new_Sorter100|7018_  = \new_Sorter100|6918_  & \new_Sorter100|6919_ ;
  assign \new_Sorter100|7019_  = \new_Sorter100|6918_  | \new_Sorter100|6919_ ;
  assign \new_Sorter100|7020_  = \new_Sorter100|6920_  & \new_Sorter100|6921_ ;
  assign \new_Sorter100|7021_  = \new_Sorter100|6920_  | \new_Sorter100|6921_ ;
  assign \new_Sorter100|7022_  = \new_Sorter100|6922_  & \new_Sorter100|6923_ ;
  assign \new_Sorter100|7023_  = \new_Sorter100|6922_  | \new_Sorter100|6923_ ;
  assign \new_Sorter100|7024_  = \new_Sorter100|6924_  & \new_Sorter100|6925_ ;
  assign \new_Sorter100|7025_  = \new_Sorter100|6924_  | \new_Sorter100|6925_ ;
  assign \new_Sorter100|7026_  = \new_Sorter100|6926_  & \new_Sorter100|6927_ ;
  assign \new_Sorter100|7027_  = \new_Sorter100|6926_  | \new_Sorter100|6927_ ;
  assign \new_Sorter100|7028_  = \new_Sorter100|6928_  & \new_Sorter100|6929_ ;
  assign \new_Sorter100|7029_  = \new_Sorter100|6928_  | \new_Sorter100|6929_ ;
  assign \new_Sorter100|7030_  = \new_Sorter100|6930_  & \new_Sorter100|6931_ ;
  assign \new_Sorter100|7031_  = \new_Sorter100|6930_  | \new_Sorter100|6931_ ;
  assign \new_Sorter100|7032_  = \new_Sorter100|6932_  & \new_Sorter100|6933_ ;
  assign \new_Sorter100|7033_  = \new_Sorter100|6932_  | \new_Sorter100|6933_ ;
  assign \new_Sorter100|7034_  = \new_Sorter100|6934_  & \new_Sorter100|6935_ ;
  assign \new_Sorter100|7035_  = \new_Sorter100|6934_  | \new_Sorter100|6935_ ;
  assign \new_Sorter100|7036_  = \new_Sorter100|6936_  & \new_Sorter100|6937_ ;
  assign \new_Sorter100|7037_  = \new_Sorter100|6936_  | \new_Sorter100|6937_ ;
  assign \new_Sorter100|7038_  = \new_Sorter100|6938_  & \new_Sorter100|6939_ ;
  assign \new_Sorter100|7039_  = \new_Sorter100|6938_  | \new_Sorter100|6939_ ;
  assign \new_Sorter100|7040_  = \new_Sorter100|6940_  & \new_Sorter100|6941_ ;
  assign \new_Sorter100|7041_  = \new_Sorter100|6940_  | \new_Sorter100|6941_ ;
  assign \new_Sorter100|7042_  = \new_Sorter100|6942_  & \new_Sorter100|6943_ ;
  assign \new_Sorter100|7043_  = \new_Sorter100|6942_  | \new_Sorter100|6943_ ;
  assign \new_Sorter100|7044_  = \new_Sorter100|6944_  & \new_Sorter100|6945_ ;
  assign \new_Sorter100|7045_  = \new_Sorter100|6944_  | \new_Sorter100|6945_ ;
  assign \new_Sorter100|7046_  = \new_Sorter100|6946_  & \new_Sorter100|6947_ ;
  assign \new_Sorter100|7047_  = \new_Sorter100|6946_  | \new_Sorter100|6947_ ;
  assign \new_Sorter100|7048_  = \new_Sorter100|6948_  & \new_Sorter100|6949_ ;
  assign \new_Sorter100|7049_  = \new_Sorter100|6948_  | \new_Sorter100|6949_ ;
  assign \new_Sorter100|7050_  = \new_Sorter100|6950_  & \new_Sorter100|6951_ ;
  assign \new_Sorter100|7051_  = \new_Sorter100|6950_  | \new_Sorter100|6951_ ;
  assign \new_Sorter100|7052_  = \new_Sorter100|6952_  & \new_Sorter100|6953_ ;
  assign \new_Sorter100|7053_  = \new_Sorter100|6952_  | \new_Sorter100|6953_ ;
  assign \new_Sorter100|7054_  = \new_Sorter100|6954_  & \new_Sorter100|6955_ ;
  assign \new_Sorter100|7055_  = \new_Sorter100|6954_  | \new_Sorter100|6955_ ;
  assign \new_Sorter100|7056_  = \new_Sorter100|6956_  & \new_Sorter100|6957_ ;
  assign \new_Sorter100|7057_  = \new_Sorter100|6956_  | \new_Sorter100|6957_ ;
  assign \new_Sorter100|7058_  = \new_Sorter100|6958_  & \new_Sorter100|6959_ ;
  assign \new_Sorter100|7059_  = \new_Sorter100|6958_  | \new_Sorter100|6959_ ;
  assign \new_Sorter100|7060_  = \new_Sorter100|6960_  & \new_Sorter100|6961_ ;
  assign \new_Sorter100|7061_  = \new_Sorter100|6960_  | \new_Sorter100|6961_ ;
  assign \new_Sorter100|7062_  = \new_Sorter100|6962_  & \new_Sorter100|6963_ ;
  assign \new_Sorter100|7063_  = \new_Sorter100|6962_  | \new_Sorter100|6963_ ;
  assign \new_Sorter100|7064_  = \new_Sorter100|6964_  & \new_Sorter100|6965_ ;
  assign \new_Sorter100|7065_  = \new_Sorter100|6964_  | \new_Sorter100|6965_ ;
  assign \new_Sorter100|7066_  = \new_Sorter100|6966_  & \new_Sorter100|6967_ ;
  assign \new_Sorter100|7067_  = \new_Sorter100|6966_  | \new_Sorter100|6967_ ;
  assign \new_Sorter100|7068_  = \new_Sorter100|6968_  & \new_Sorter100|6969_ ;
  assign \new_Sorter100|7069_  = \new_Sorter100|6968_  | \new_Sorter100|6969_ ;
  assign \new_Sorter100|7070_  = \new_Sorter100|6970_  & \new_Sorter100|6971_ ;
  assign \new_Sorter100|7071_  = \new_Sorter100|6970_  | \new_Sorter100|6971_ ;
  assign \new_Sorter100|7072_  = \new_Sorter100|6972_  & \new_Sorter100|6973_ ;
  assign \new_Sorter100|7073_  = \new_Sorter100|6972_  | \new_Sorter100|6973_ ;
  assign \new_Sorter100|7074_  = \new_Sorter100|6974_  & \new_Sorter100|6975_ ;
  assign \new_Sorter100|7075_  = \new_Sorter100|6974_  | \new_Sorter100|6975_ ;
  assign \new_Sorter100|7076_  = \new_Sorter100|6976_  & \new_Sorter100|6977_ ;
  assign \new_Sorter100|7077_  = \new_Sorter100|6976_  | \new_Sorter100|6977_ ;
  assign \new_Sorter100|7078_  = \new_Sorter100|6978_  & \new_Sorter100|6979_ ;
  assign \new_Sorter100|7079_  = \new_Sorter100|6978_  | \new_Sorter100|6979_ ;
  assign \new_Sorter100|7080_  = \new_Sorter100|6980_  & \new_Sorter100|6981_ ;
  assign \new_Sorter100|7081_  = \new_Sorter100|6980_  | \new_Sorter100|6981_ ;
  assign \new_Sorter100|7082_  = \new_Sorter100|6982_  & \new_Sorter100|6983_ ;
  assign \new_Sorter100|7083_  = \new_Sorter100|6982_  | \new_Sorter100|6983_ ;
  assign \new_Sorter100|7084_  = \new_Sorter100|6984_  & \new_Sorter100|6985_ ;
  assign \new_Sorter100|7085_  = \new_Sorter100|6984_  | \new_Sorter100|6985_ ;
  assign \new_Sorter100|7086_  = \new_Sorter100|6986_  & \new_Sorter100|6987_ ;
  assign \new_Sorter100|7087_  = \new_Sorter100|6986_  | \new_Sorter100|6987_ ;
  assign \new_Sorter100|7088_  = \new_Sorter100|6988_  & \new_Sorter100|6989_ ;
  assign \new_Sorter100|7089_  = \new_Sorter100|6988_  | \new_Sorter100|6989_ ;
  assign \new_Sorter100|7090_  = \new_Sorter100|6990_  & \new_Sorter100|6991_ ;
  assign \new_Sorter100|7091_  = \new_Sorter100|6990_  | \new_Sorter100|6991_ ;
  assign \new_Sorter100|7092_  = \new_Sorter100|6992_  & \new_Sorter100|6993_ ;
  assign \new_Sorter100|7093_  = \new_Sorter100|6992_  | \new_Sorter100|6993_ ;
  assign \new_Sorter100|7094_  = \new_Sorter100|6994_  & \new_Sorter100|6995_ ;
  assign \new_Sorter100|7095_  = \new_Sorter100|6994_  | \new_Sorter100|6995_ ;
  assign \new_Sorter100|7096_  = \new_Sorter100|6996_  & \new_Sorter100|6997_ ;
  assign \new_Sorter100|7097_  = \new_Sorter100|6996_  | \new_Sorter100|6997_ ;
  assign \new_Sorter100|7098_  = \new_Sorter100|6998_  & \new_Sorter100|6999_ ;
  assign \new_Sorter100|7099_  = \new_Sorter100|6998_  | \new_Sorter100|6999_ ;
  assign \new_Sorter100|7100_  = \new_Sorter100|7000_ ;
  assign \new_Sorter100|7199_  = \new_Sorter100|7099_ ;
  assign \new_Sorter100|7101_  = \new_Sorter100|7001_  & \new_Sorter100|7002_ ;
  assign \new_Sorter100|7102_  = \new_Sorter100|7001_  | \new_Sorter100|7002_ ;
  assign \new_Sorter100|7103_  = \new_Sorter100|7003_  & \new_Sorter100|7004_ ;
  assign \new_Sorter100|7104_  = \new_Sorter100|7003_  | \new_Sorter100|7004_ ;
  assign \new_Sorter100|7105_  = \new_Sorter100|7005_  & \new_Sorter100|7006_ ;
  assign \new_Sorter100|7106_  = \new_Sorter100|7005_  | \new_Sorter100|7006_ ;
  assign \new_Sorter100|7107_  = \new_Sorter100|7007_  & \new_Sorter100|7008_ ;
  assign \new_Sorter100|7108_  = \new_Sorter100|7007_  | \new_Sorter100|7008_ ;
  assign \new_Sorter100|7109_  = \new_Sorter100|7009_  & \new_Sorter100|7010_ ;
  assign \new_Sorter100|7110_  = \new_Sorter100|7009_  | \new_Sorter100|7010_ ;
  assign \new_Sorter100|7111_  = \new_Sorter100|7011_  & \new_Sorter100|7012_ ;
  assign \new_Sorter100|7112_  = \new_Sorter100|7011_  | \new_Sorter100|7012_ ;
  assign \new_Sorter100|7113_  = \new_Sorter100|7013_  & \new_Sorter100|7014_ ;
  assign \new_Sorter100|7114_  = \new_Sorter100|7013_  | \new_Sorter100|7014_ ;
  assign \new_Sorter100|7115_  = \new_Sorter100|7015_  & \new_Sorter100|7016_ ;
  assign \new_Sorter100|7116_  = \new_Sorter100|7015_  | \new_Sorter100|7016_ ;
  assign \new_Sorter100|7117_  = \new_Sorter100|7017_  & \new_Sorter100|7018_ ;
  assign \new_Sorter100|7118_  = \new_Sorter100|7017_  | \new_Sorter100|7018_ ;
  assign \new_Sorter100|7119_  = \new_Sorter100|7019_  & \new_Sorter100|7020_ ;
  assign \new_Sorter100|7120_  = \new_Sorter100|7019_  | \new_Sorter100|7020_ ;
  assign \new_Sorter100|7121_  = \new_Sorter100|7021_  & \new_Sorter100|7022_ ;
  assign \new_Sorter100|7122_  = \new_Sorter100|7021_  | \new_Sorter100|7022_ ;
  assign \new_Sorter100|7123_  = \new_Sorter100|7023_  & \new_Sorter100|7024_ ;
  assign \new_Sorter100|7124_  = \new_Sorter100|7023_  | \new_Sorter100|7024_ ;
  assign \new_Sorter100|7125_  = \new_Sorter100|7025_  & \new_Sorter100|7026_ ;
  assign \new_Sorter100|7126_  = \new_Sorter100|7025_  | \new_Sorter100|7026_ ;
  assign \new_Sorter100|7127_  = \new_Sorter100|7027_  & \new_Sorter100|7028_ ;
  assign \new_Sorter100|7128_  = \new_Sorter100|7027_  | \new_Sorter100|7028_ ;
  assign \new_Sorter100|7129_  = \new_Sorter100|7029_  & \new_Sorter100|7030_ ;
  assign \new_Sorter100|7130_  = \new_Sorter100|7029_  | \new_Sorter100|7030_ ;
  assign \new_Sorter100|7131_  = \new_Sorter100|7031_  & \new_Sorter100|7032_ ;
  assign \new_Sorter100|7132_  = \new_Sorter100|7031_  | \new_Sorter100|7032_ ;
  assign \new_Sorter100|7133_  = \new_Sorter100|7033_  & \new_Sorter100|7034_ ;
  assign \new_Sorter100|7134_  = \new_Sorter100|7033_  | \new_Sorter100|7034_ ;
  assign \new_Sorter100|7135_  = \new_Sorter100|7035_  & \new_Sorter100|7036_ ;
  assign \new_Sorter100|7136_  = \new_Sorter100|7035_  | \new_Sorter100|7036_ ;
  assign \new_Sorter100|7137_  = \new_Sorter100|7037_  & \new_Sorter100|7038_ ;
  assign \new_Sorter100|7138_  = \new_Sorter100|7037_  | \new_Sorter100|7038_ ;
  assign \new_Sorter100|7139_  = \new_Sorter100|7039_  & \new_Sorter100|7040_ ;
  assign \new_Sorter100|7140_  = \new_Sorter100|7039_  | \new_Sorter100|7040_ ;
  assign \new_Sorter100|7141_  = \new_Sorter100|7041_  & \new_Sorter100|7042_ ;
  assign \new_Sorter100|7142_  = \new_Sorter100|7041_  | \new_Sorter100|7042_ ;
  assign \new_Sorter100|7143_  = \new_Sorter100|7043_  & \new_Sorter100|7044_ ;
  assign \new_Sorter100|7144_  = \new_Sorter100|7043_  | \new_Sorter100|7044_ ;
  assign \new_Sorter100|7145_  = \new_Sorter100|7045_  & \new_Sorter100|7046_ ;
  assign \new_Sorter100|7146_  = \new_Sorter100|7045_  | \new_Sorter100|7046_ ;
  assign \new_Sorter100|7147_  = \new_Sorter100|7047_  & \new_Sorter100|7048_ ;
  assign \new_Sorter100|7148_  = \new_Sorter100|7047_  | \new_Sorter100|7048_ ;
  assign \new_Sorter100|7149_  = \new_Sorter100|7049_  & \new_Sorter100|7050_ ;
  assign \new_Sorter100|7150_  = \new_Sorter100|7049_  | \new_Sorter100|7050_ ;
  assign \new_Sorter100|7151_  = \new_Sorter100|7051_  & \new_Sorter100|7052_ ;
  assign \new_Sorter100|7152_  = \new_Sorter100|7051_  | \new_Sorter100|7052_ ;
  assign \new_Sorter100|7153_  = \new_Sorter100|7053_  & \new_Sorter100|7054_ ;
  assign \new_Sorter100|7154_  = \new_Sorter100|7053_  | \new_Sorter100|7054_ ;
  assign \new_Sorter100|7155_  = \new_Sorter100|7055_  & \new_Sorter100|7056_ ;
  assign \new_Sorter100|7156_  = \new_Sorter100|7055_  | \new_Sorter100|7056_ ;
  assign \new_Sorter100|7157_  = \new_Sorter100|7057_  & \new_Sorter100|7058_ ;
  assign \new_Sorter100|7158_  = \new_Sorter100|7057_  | \new_Sorter100|7058_ ;
  assign \new_Sorter100|7159_  = \new_Sorter100|7059_  & \new_Sorter100|7060_ ;
  assign \new_Sorter100|7160_  = \new_Sorter100|7059_  | \new_Sorter100|7060_ ;
  assign \new_Sorter100|7161_  = \new_Sorter100|7061_  & \new_Sorter100|7062_ ;
  assign \new_Sorter100|7162_  = \new_Sorter100|7061_  | \new_Sorter100|7062_ ;
  assign \new_Sorter100|7163_  = \new_Sorter100|7063_  & \new_Sorter100|7064_ ;
  assign \new_Sorter100|7164_  = \new_Sorter100|7063_  | \new_Sorter100|7064_ ;
  assign \new_Sorter100|7165_  = \new_Sorter100|7065_  & \new_Sorter100|7066_ ;
  assign \new_Sorter100|7166_  = \new_Sorter100|7065_  | \new_Sorter100|7066_ ;
  assign \new_Sorter100|7167_  = \new_Sorter100|7067_  & \new_Sorter100|7068_ ;
  assign \new_Sorter100|7168_  = \new_Sorter100|7067_  | \new_Sorter100|7068_ ;
  assign \new_Sorter100|7169_  = \new_Sorter100|7069_  & \new_Sorter100|7070_ ;
  assign \new_Sorter100|7170_  = \new_Sorter100|7069_  | \new_Sorter100|7070_ ;
  assign \new_Sorter100|7171_  = \new_Sorter100|7071_  & \new_Sorter100|7072_ ;
  assign \new_Sorter100|7172_  = \new_Sorter100|7071_  | \new_Sorter100|7072_ ;
  assign \new_Sorter100|7173_  = \new_Sorter100|7073_  & \new_Sorter100|7074_ ;
  assign \new_Sorter100|7174_  = \new_Sorter100|7073_  | \new_Sorter100|7074_ ;
  assign \new_Sorter100|7175_  = \new_Sorter100|7075_  & \new_Sorter100|7076_ ;
  assign \new_Sorter100|7176_  = \new_Sorter100|7075_  | \new_Sorter100|7076_ ;
  assign \new_Sorter100|7177_  = \new_Sorter100|7077_  & \new_Sorter100|7078_ ;
  assign \new_Sorter100|7178_  = \new_Sorter100|7077_  | \new_Sorter100|7078_ ;
  assign \new_Sorter100|7179_  = \new_Sorter100|7079_  & \new_Sorter100|7080_ ;
  assign \new_Sorter100|7180_  = \new_Sorter100|7079_  | \new_Sorter100|7080_ ;
  assign \new_Sorter100|7181_  = \new_Sorter100|7081_  & \new_Sorter100|7082_ ;
  assign \new_Sorter100|7182_  = \new_Sorter100|7081_  | \new_Sorter100|7082_ ;
  assign \new_Sorter100|7183_  = \new_Sorter100|7083_  & \new_Sorter100|7084_ ;
  assign \new_Sorter100|7184_  = \new_Sorter100|7083_  | \new_Sorter100|7084_ ;
  assign \new_Sorter100|7185_  = \new_Sorter100|7085_  & \new_Sorter100|7086_ ;
  assign \new_Sorter100|7186_  = \new_Sorter100|7085_  | \new_Sorter100|7086_ ;
  assign \new_Sorter100|7187_  = \new_Sorter100|7087_  & \new_Sorter100|7088_ ;
  assign \new_Sorter100|7188_  = \new_Sorter100|7087_  | \new_Sorter100|7088_ ;
  assign \new_Sorter100|7189_  = \new_Sorter100|7089_  & \new_Sorter100|7090_ ;
  assign \new_Sorter100|7190_  = \new_Sorter100|7089_  | \new_Sorter100|7090_ ;
  assign \new_Sorter100|7191_  = \new_Sorter100|7091_  & \new_Sorter100|7092_ ;
  assign \new_Sorter100|7192_  = \new_Sorter100|7091_  | \new_Sorter100|7092_ ;
  assign \new_Sorter100|7193_  = \new_Sorter100|7093_  & \new_Sorter100|7094_ ;
  assign \new_Sorter100|7194_  = \new_Sorter100|7093_  | \new_Sorter100|7094_ ;
  assign \new_Sorter100|7195_  = \new_Sorter100|7095_  & \new_Sorter100|7096_ ;
  assign \new_Sorter100|7196_  = \new_Sorter100|7095_  | \new_Sorter100|7096_ ;
  assign \new_Sorter100|7197_  = \new_Sorter100|7097_  & \new_Sorter100|7098_ ;
  assign \new_Sorter100|7198_  = \new_Sorter100|7097_  | \new_Sorter100|7098_ ;
  assign \new_Sorter100|7200_  = \new_Sorter100|7100_  & \new_Sorter100|7101_ ;
  assign \new_Sorter100|7201_  = \new_Sorter100|7100_  | \new_Sorter100|7101_ ;
  assign \new_Sorter100|7202_  = \new_Sorter100|7102_  & \new_Sorter100|7103_ ;
  assign \new_Sorter100|7203_  = \new_Sorter100|7102_  | \new_Sorter100|7103_ ;
  assign \new_Sorter100|7204_  = \new_Sorter100|7104_  & \new_Sorter100|7105_ ;
  assign \new_Sorter100|7205_  = \new_Sorter100|7104_  | \new_Sorter100|7105_ ;
  assign \new_Sorter100|7206_  = \new_Sorter100|7106_  & \new_Sorter100|7107_ ;
  assign \new_Sorter100|7207_  = \new_Sorter100|7106_  | \new_Sorter100|7107_ ;
  assign \new_Sorter100|7208_  = \new_Sorter100|7108_  & \new_Sorter100|7109_ ;
  assign \new_Sorter100|7209_  = \new_Sorter100|7108_  | \new_Sorter100|7109_ ;
  assign \new_Sorter100|7210_  = \new_Sorter100|7110_  & \new_Sorter100|7111_ ;
  assign \new_Sorter100|7211_  = \new_Sorter100|7110_  | \new_Sorter100|7111_ ;
  assign \new_Sorter100|7212_  = \new_Sorter100|7112_  & \new_Sorter100|7113_ ;
  assign \new_Sorter100|7213_  = \new_Sorter100|7112_  | \new_Sorter100|7113_ ;
  assign \new_Sorter100|7214_  = \new_Sorter100|7114_  & \new_Sorter100|7115_ ;
  assign \new_Sorter100|7215_  = \new_Sorter100|7114_  | \new_Sorter100|7115_ ;
  assign \new_Sorter100|7216_  = \new_Sorter100|7116_  & \new_Sorter100|7117_ ;
  assign \new_Sorter100|7217_  = \new_Sorter100|7116_  | \new_Sorter100|7117_ ;
  assign \new_Sorter100|7218_  = \new_Sorter100|7118_  & \new_Sorter100|7119_ ;
  assign \new_Sorter100|7219_  = \new_Sorter100|7118_  | \new_Sorter100|7119_ ;
  assign \new_Sorter100|7220_  = \new_Sorter100|7120_  & \new_Sorter100|7121_ ;
  assign \new_Sorter100|7221_  = \new_Sorter100|7120_  | \new_Sorter100|7121_ ;
  assign \new_Sorter100|7222_  = \new_Sorter100|7122_  & \new_Sorter100|7123_ ;
  assign \new_Sorter100|7223_  = \new_Sorter100|7122_  | \new_Sorter100|7123_ ;
  assign \new_Sorter100|7224_  = \new_Sorter100|7124_  & \new_Sorter100|7125_ ;
  assign \new_Sorter100|7225_  = \new_Sorter100|7124_  | \new_Sorter100|7125_ ;
  assign \new_Sorter100|7226_  = \new_Sorter100|7126_  & \new_Sorter100|7127_ ;
  assign \new_Sorter100|7227_  = \new_Sorter100|7126_  | \new_Sorter100|7127_ ;
  assign \new_Sorter100|7228_  = \new_Sorter100|7128_  & \new_Sorter100|7129_ ;
  assign \new_Sorter100|7229_  = \new_Sorter100|7128_  | \new_Sorter100|7129_ ;
  assign \new_Sorter100|7230_  = \new_Sorter100|7130_  & \new_Sorter100|7131_ ;
  assign \new_Sorter100|7231_  = \new_Sorter100|7130_  | \new_Sorter100|7131_ ;
  assign \new_Sorter100|7232_  = \new_Sorter100|7132_  & \new_Sorter100|7133_ ;
  assign \new_Sorter100|7233_  = \new_Sorter100|7132_  | \new_Sorter100|7133_ ;
  assign \new_Sorter100|7234_  = \new_Sorter100|7134_  & \new_Sorter100|7135_ ;
  assign \new_Sorter100|7235_  = \new_Sorter100|7134_  | \new_Sorter100|7135_ ;
  assign \new_Sorter100|7236_  = \new_Sorter100|7136_  & \new_Sorter100|7137_ ;
  assign \new_Sorter100|7237_  = \new_Sorter100|7136_  | \new_Sorter100|7137_ ;
  assign \new_Sorter100|7238_  = \new_Sorter100|7138_  & \new_Sorter100|7139_ ;
  assign \new_Sorter100|7239_  = \new_Sorter100|7138_  | \new_Sorter100|7139_ ;
  assign \new_Sorter100|7240_  = \new_Sorter100|7140_  & \new_Sorter100|7141_ ;
  assign \new_Sorter100|7241_  = \new_Sorter100|7140_  | \new_Sorter100|7141_ ;
  assign \new_Sorter100|7242_  = \new_Sorter100|7142_  & \new_Sorter100|7143_ ;
  assign \new_Sorter100|7243_  = \new_Sorter100|7142_  | \new_Sorter100|7143_ ;
  assign \new_Sorter100|7244_  = \new_Sorter100|7144_  & \new_Sorter100|7145_ ;
  assign \new_Sorter100|7245_  = \new_Sorter100|7144_  | \new_Sorter100|7145_ ;
  assign \new_Sorter100|7246_  = \new_Sorter100|7146_  & \new_Sorter100|7147_ ;
  assign \new_Sorter100|7247_  = \new_Sorter100|7146_  | \new_Sorter100|7147_ ;
  assign \new_Sorter100|7248_  = \new_Sorter100|7148_  & \new_Sorter100|7149_ ;
  assign \new_Sorter100|7249_  = \new_Sorter100|7148_  | \new_Sorter100|7149_ ;
  assign \new_Sorter100|7250_  = \new_Sorter100|7150_  & \new_Sorter100|7151_ ;
  assign \new_Sorter100|7251_  = \new_Sorter100|7150_  | \new_Sorter100|7151_ ;
  assign \new_Sorter100|7252_  = \new_Sorter100|7152_  & \new_Sorter100|7153_ ;
  assign \new_Sorter100|7253_  = \new_Sorter100|7152_  | \new_Sorter100|7153_ ;
  assign \new_Sorter100|7254_  = \new_Sorter100|7154_  & \new_Sorter100|7155_ ;
  assign \new_Sorter100|7255_  = \new_Sorter100|7154_  | \new_Sorter100|7155_ ;
  assign \new_Sorter100|7256_  = \new_Sorter100|7156_  & \new_Sorter100|7157_ ;
  assign \new_Sorter100|7257_  = \new_Sorter100|7156_  | \new_Sorter100|7157_ ;
  assign \new_Sorter100|7258_  = \new_Sorter100|7158_  & \new_Sorter100|7159_ ;
  assign \new_Sorter100|7259_  = \new_Sorter100|7158_  | \new_Sorter100|7159_ ;
  assign \new_Sorter100|7260_  = \new_Sorter100|7160_  & \new_Sorter100|7161_ ;
  assign \new_Sorter100|7261_  = \new_Sorter100|7160_  | \new_Sorter100|7161_ ;
  assign \new_Sorter100|7262_  = \new_Sorter100|7162_  & \new_Sorter100|7163_ ;
  assign \new_Sorter100|7263_  = \new_Sorter100|7162_  | \new_Sorter100|7163_ ;
  assign \new_Sorter100|7264_  = \new_Sorter100|7164_  & \new_Sorter100|7165_ ;
  assign \new_Sorter100|7265_  = \new_Sorter100|7164_  | \new_Sorter100|7165_ ;
  assign \new_Sorter100|7266_  = \new_Sorter100|7166_  & \new_Sorter100|7167_ ;
  assign \new_Sorter100|7267_  = \new_Sorter100|7166_  | \new_Sorter100|7167_ ;
  assign \new_Sorter100|7268_  = \new_Sorter100|7168_  & \new_Sorter100|7169_ ;
  assign \new_Sorter100|7269_  = \new_Sorter100|7168_  | \new_Sorter100|7169_ ;
  assign \new_Sorter100|7270_  = \new_Sorter100|7170_  & \new_Sorter100|7171_ ;
  assign \new_Sorter100|7271_  = \new_Sorter100|7170_  | \new_Sorter100|7171_ ;
  assign \new_Sorter100|7272_  = \new_Sorter100|7172_  & \new_Sorter100|7173_ ;
  assign \new_Sorter100|7273_  = \new_Sorter100|7172_  | \new_Sorter100|7173_ ;
  assign \new_Sorter100|7274_  = \new_Sorter100|7174_  & \new_Sorter100|7175_ ;
  assign \new_Sorter100|7275_  = \new_Sorter100|7174_  | \new_Sorter100|7175_ ;
  assign \new_Sorter100|7276_  = \new_Sorter100|7176_  & \new_Sorter100|7177_ ;
  assign \new_Sorter100|7277_  = \new_Sorter100|7176_  | \new_Sorter100|7177_ ;
  assign \new_Sorter100|7278_  = \new_Sorter100|7178_  & \new_Sorter100|7179_ ;
  assign \new_Sorter100|7279_  = \new_Sorter100|7178_  | \new_Sorter100|7179_ ;
  assign \new_Sorter100|7280_  = \new_Sorter100|7180_  & \new_Sorter100|7181_ ;
  assign \new_Sorter100|7281_  = \new_Sorter100|7180_  | \new_Sorter100|7181_ ;
  assign \new_Sorter100|7282_  = \new_Sorter100|7182_  & \new_Sorter100|7183_ ;
  assign \new_Sorter100|7283_  = \new_Sorter100|7182_  | \new_Sorter100|7183_ ;
  assign \new_Sorter100|7284_  = \new_Sorter100|7184_  & \new_Sorter100|7185_ ;
  assign \new_Sorter100|7285_  = \new_Sorter100|7184_  | \new_Sorter100|7185_ ;
  assign \new_Sorter100|7286_  = \new_Sorter100|7186_  & \new_Sorter100|7187_ ;
  assign \new_Sorter100|7287_  = \new_Sorter100|7186_  | \new_Sorter100|7187_ ;
  assign \new_Sorter100|7288_  = \new_Sorter100|7188_  & \new_Sorter100|7189_ ;
  assign \new_Sorter100|7289_  = \new_Sorter100|7188_  | \new_Sorter100|7189_ ;
  assign \new_Sorter100|7290_  = \new_Sorter100|7190_  & \new_Sorter100|7191_ ;
  assign \new_Sorter100|7291_  = \new_Sorter100|7190_  | \new_Sorter100|7191_ ;
  assign \new_Sorter100|7292_  = \new_Sorter100|7192_  & \new_Sorter100|7193_ ;
  assign \new_Sorter100|7293_  = \new_Sorter100|7192_  | \new_Sorter100|7193_ ;
  assign \new_Sorter100|7294_  = \new_Sorter100|7194_  & \new_Sorter100|7195_ ;
  assign \new_Sorter100|7295_  = \new_Sorter100|7194_  | \new_Sorter100|7195_ ;
  assign \new_Sorter100|7296_  = \new_Sorter100|7196_  & \new_Sorter100|7197_ ;
  assign \new_Sorter100|7297_  = \new_Sorter100|7196_  | \new_Sorter100|7197_ ;
  assign \new_Sorter100|7298_  = \new_Sorter100|7198_  & \new_Sorter100|7199_ ;
  assign \new_Sorter100|7299_  = \new_Sorter100|7198_  | \new_Sorter100|7199_ ;
  assign \new_Sorter100|7300_  = \new_Sorter100|7200_ ;
  assign \new_Sorter100|7399_  = \new_Sorter100|7299_ ;
  assign \new_Sorter100|7301_  = \new_Sorter100|7201_  & \new_Sorter100|7202_ ;
  assign \new_Sorter100|7302_  = \new_Sorter100|7201_  | \new_Sorter100|7202_ ;
  assign \new_Sorter100|7303_  = \new_Sorter100|7203_  & \new_Sorter100|7204_ ;
  assign \new_Sorter100|7304_  = \new_Sorter100|7203_  | \new_Sorter100|7204_ ;
  assign \new_Sorter100|7305_  = \new_Sorter100|7205_  & \new_Sorter100|7206_ ;
  assign \new_Sorter100|7306_  = \new_Sorter100|7205_  | \new_Sorter100|7206_ ;
  assign \new_Sorter100|7307_  = \new_Sorter100|7207_  & \new_Sorter100|7208_ ;
  assign \new_Sorter100|7308_  = \new_Sorter100|7207_  | \new_Sorter100|7208_ ;
  assign \new_Sorter100|7309_  = \new_Sorter100|7209_  & \new_Sorter100|7210_ ;
  assign \new_Sorter100|7310_  = \new_Sorter100|7209_  | \new_Sorter100|7210_ ;
  assign \new_Sorter100|7311_  = \new_Sorter100|7211_  & \new_Sorter100|7212_ ;
  assign \new_Sorter100|7312_  = \new_Sorter100|7211_  | \new_Sorter100|7212_ ;
  assign \new_Sorter100|7313_  = \new_Sorter100|7213_  & \new_Sorter100|7214_ ;
  assign \new_Sorter100|7314_  = \new_Sorter100|7213_  | \new_Sorter100|7214_ ;
  assign \new_Sorter100|7315_  = \new_Sorter100|7215_  & \new_Sorter100|7216_ ;
  assign \new_Sorter100|7316_  = \new_Sorter100|7215_  | \new_Sorter100|7216_ ;
  assign \new_Sorter100|7317_  = \new_Sorter100|7217_  & \new_Sorter100|7218_ ;
  assign \new_Sorter100|7318_  = \new_Sorter100|7217_  | \new_Sorter100|7218_ ;
  assign \new_Sorter100|7319_  = \new_Sorter100|7219_  & \new_Sorter100|7220_ ;
  assign \new_Sorter100|7320_  = \new_Sorter100|7219_  | \new_Sorter100|7220_ ;
  assign \new_Sorter100|7321_  = \new_Sorter100|7221_  & \new_Sorter100|7222_ ;
  assign \new_Sorter100|7322_  = \new_Sorter100|7221_  | \new_Sorter100|7222_ ;
  assign \new_Sorter100|7323_  = \new_Sorter100|7223_  & \new_Sorter100|7224_ ;
  assign \new_Sorter100|7324_  = \new_Sorter100|7223_  | \new_Sorter100|7224_ ;
  assign \new_Sorter100|7325_  = \new_Sorter100|7225_  & \new_Sorter100|7226_ ;
  assign \new_Sorter100|7326_  = \new_Sorter100|7225_  | \new_Sorter100|7226_ ;
  assign \new_Sorter100|7327_  = \new_Sorter100|7227_  & \new_Sorter100|7228_ ;
  assign \new_Sorter100|7328_  = \new_Sorter100|7227_  | \new_Sorter100|7228_ ;
  assign \new_Sorter100|7329_  = \new_Sorter100|7229_  & \new_Sorter100|7230_ ;
  assign \new_Sorter100|7330_  = \new_Sorter100|7229_  | \new_Sorter100|7230_ ;
  assign \new_Sorter100|7331_  = \new_Sorter100|7231_  & \new_Sorter100|7232_ ;
  assign \new_Sorter100|7332_  = \new_Sorter100|7231_  | \new_Sorter100|7232_ ;
  assign \new_Sorter100|7333_  = \new_Sorter100|7233_  & \new_Sorter100|7234_ ;
  assign \new_Sorter100|7334_  = \new_Sorter100|7233_  | \new_Sorter100|7234_ ;
  assign \new_Sorter100|7335_  = \new_Sorter100|7235_  & \new_Sorter100|7236_ ;
  assign \new_Sorter100|7336_  = \new_Sorter100|7235_  | \new_Sorter100|7236_ ;
  assign \new_Sorter100|7337_  = \new_Sorter100|7237_  & \new_Sorter100|7238_ ;
  assign \new_Sorter100|7338_  = \new_Sorter100|7237_  | \new_Sorter100|7238_ ;
  assign \new_Sorter100|7339_  = \new_Sorter100|7239_  & \new_Sorter100|7240_ ;
  assign \new_Sorter100|7340_  = \new_Sorter100|7239_  | \new_Sorter100|7240_ ;
  assign \new_Sorter100|7341_  = \new_Sorter100|7241_  & \new_Sorter100|7242_ ;
  assign \new_Sorter100|7342_  = \new_Sorter100|7241_  | \new_Sorter100|7242_ ;
  assign \new_Sorter100|7343_  = \new_Sorter100|7243_  & \new_Sorter100|7244_ ;
  assign \new_Sorter100|7344_  = \new_Sorter100|7243_  | \new_Sorter100|7244_ ;
  assign \new_Sorter100|7345_  = \new_Sorter100|7245_  & \new_Sorter100|7246_ ;
  assign \new_Sorter100|7346_  = \new_Sorter100|7245_  | \new_Sorter100|7246_ ;
  assign \new_Sorter100|7347_  = \new_Sorter100|7247_  & \new_Sorter100|7248_ ;
  assign \new_Sorter100|7348_  = \new_Sorter100|7247_  | \new_Sorter100|7248_ ;
  assign \new_Sorter100|7349_  = \new_Sorter100|7249_  & \new_Sorter100|7250_ ;
  assign \new_Sorter100|7350_  = \new_Sorter100|7249_  | \new_Sorter100|7250_ ;
  assign \new_Sorter100|7351_  = \new_Sorter100|7251_  & \new_Sorter100|7252_ ;
  assign \new_Sorter100|7352_  = \new_Sorter100|7251_  | \new_Sorter100|7252_ ;
  assign \new_Sorter100|7353_  = \new_Sorter100|7253_  & \new_Sorter100|7254_ ;
  assign \new_Sorter100|7354_  = \new_Sorter100|7253_  | \new_Sorter100|7254_ ;
  assign \new_Sorter100|7355_  = \new_Sorter100|7255_  & \new_Sorter100|7256_ ;
  assign \new_Sorter100|7356_  = \new_Sorter100|7255_  | \new_Sorter100|7256_ ;
  assign \new_Sorter100|7357_  = \new_Sorter100|7257_  & \new_Sorter100|7258_ ;
  assign \new_Sorter100|7358_  = \new_Sorter100|7257_  | \new_Sorter100|7258_ ;
  assign \new_Sorter100|7359_  = \new_Sorter100|7259_  & \new_Sorter100|7260_ ;
  assign \new_Sorter100|7360_  = \new_Sorter100|7259_  | \new_Sorter100|7260_ ;
  assign \new_Sorter100|7361_  = \new_Sorter100|7261_  & \new_Sorter100|7262_ ;
  assign \new_Sorter100|7362_  = \new_Sorter100|7261_  | \new_Sorter100|7262_ ;
  assign \new_Sorter100|7363_  = \new_Sorter100|7263_  & \new_Sorter100|7264_ ;
  assign \new_Sorter100|7364_  = \new_Sorter100|7263_  | \new_Sorter100|7264_ ;
  assign \new_Sorter100|7365_  = \new_Sorter100|7265_  & \new_Sorter100|7266_ ;
  assign \new_Sorter100|7366_  = \new_Sorter100|7265_  | \new_Sorter100|7266_ ;
  assign \new_Sorter100|7367_  = \new_Sorter100|7267_  & \new_Sorter100|7268_ ;
  assign \new_Sorter100|7368_  = \new_Sorter100|7267_  | \new_Sorter100|7268_ ;
  assign \new_Sorter100|7369_  = \new_Sorter100|7269_  & \new_Sorter100|7270_ ;
  assign \new_Sorter100|7370_  = \new_Sorter100|7269_  | \new_Sorter100|7270_ ;
  assign \new_Sorter100|7371_  = \new_Sorter100|7271_  & \new_Sorter100|7272_ ;
  assign \new_Sorter100|7372_  = \new_Sorter100|7271_  | \new_Sorter100|7272_ ;
  assign \new_Sorter100|7373_  = \new_Sorter100|7273_  & \new_Sorter100|7274_ ;
  assign \new_Sorter100|7374_  = \new_Sorter100|7273_  | \new_Sorter100|7274_ ;
  assign \new_Sorter100|7375_  = \new_Sorter100|7275_  & \new_Sorter100|7276_ ;
  assign \new_Sorter100|7376_  = \new_Sorter100|7275_  | \new_Sorter100|7276_ ;
  assign \new_Sorter100|7377_  = \new_Sorter100|7277_  & \new_Sorter100|7278_ ;
  assign \new_Sorter100|7378_  = \new_Sorter100|7277_  | \new_Sorter100|7278_ ;
  assign \new_Sorter100|7379_  = \new_Sorter100|7279_  & \new_Sorter100|7280_ ;
  assign \new_Sorter100|7380_  = \new_Sorter100|7279_  | \new_Sorter100|7280_ ;
  assign \new_Sorter100|7381_  = \new_Sorter100|7281_  & \new_Sorter100|7282_ ;
  assign \new_Sorter100|7382_  = \new_Sorter100|7281_  | \new_Sorter100|7282_ ;
  assign \new_Sorter100|7383_  = \new_Sorter100|7283_  & \new_Sorter100|7284_ ;
  assign \new_Sorter100|7384_  = \new_Sorter100|7283_  | \new_Sorter100|7284_ ;
  assign \new_Sorter100|7385_  = \new_Sorter100|7285_  & \new_Sorter100|7286_ ;
  assign \new_Sorter100|7386_  = \new_Sorter100|7285_  | \new_Sorter100|7286_ ;
  assign \new_Sorter100|7387_  = \new_Sorter100|7287_  & \new_Sorter100|7288_ ;
  assign \new_Sorter100|7388_  = \new_Sorter100|7287_  | \new_Sorter100|7288_ ;
  assign \new_Sorter100|7389_  = \new_Sorter100|7289_  & \new_Sorter100|7290_ ;
  assign \new_Sorter100|7390_  = \new_Sorter100|7289_  | \new_Sorter100|7290_ ;
  assign \new_Sorter100|7391_  = \new_Sorter100|7291_  & \new_Sorter100|7292_ ;
  assign \new_Sorter100|7392_  = \new_Sorter100|7291_  | \new_Sorter100|7292_ ;
  assign \new_Sorter100|7393_  = \new_Sorter100|7293_  & \new_Sorter100|7294_ ;
  assign \new_Sorter100|7394_  = \new_Sorter100|7293_  | \new_Sorter100|7294_ ;
  assign \new_Sorter100|7395_  = \new_Sorter100|7295_  & \new_Sorter100|7296_ ;
  assign \new_Sorter100|7396_  = \new_Sorter100|7295_  | \new_Sorter100|7296_ ;
  assign \new_Sorter100|7397_  = \new_Sorter100|7297_  & \new_Sorter100|7298_ ;
  assign \new_Sorter100|7398_  = \new_Sorter100|7297_  | \new_Sorter100|7298_ ;
  assign \new_Sorter100|7400_  = \new_Sorter100|7300_  & \new_Sorter100|7301_ ;
  assign \new_Sorter100|7401_  = \new_Sorter100|7300_  | \new_Sorter100|7301_ ;
  assign \new_Sorter100|7402_  = \new_Sorter100|7302_  & \new_Sorter100|7303_ ;
  assign \new_Sorter100|7403_  = \new_Sorter100|7302_  | \new_Sorter100|7303_ ;
  assign \new_Sorter100|7404_  = \new_Sorter100|7304_  & \new_Sorter100|7305_ ;
  assign \new_Sorter100|7405_  = \new_Sorter100|7304_  | \new_Sorter100|7305_ ;
  assign \new_Sorter100|7406_  = \new_Sorter100|7306_  & \new_Sorter100|7307_ ;
  assign \new_Sorter100|7407_  = \new_Sorter100|7306_  | \new_Sorter100|7307_ ;
  assign \new_Sorter100|7408_  = \new_Sorter100|7308_  & \new_Sorter100|7309_ ;
  assign \new_Sorter100|7409_  = \new_Sorter100|7308_  | \new_Sorter100|7309_ ;
  assign \new_Sorter100|7410_  = \new_Sorter100|7310_  & \new_Sorter100|7311_ ;
  assign \new_Sorter100|7411_  = \new_Sorter100|7310_  | \new_Sorter100|7311_ ;
  assign \new_Sorter100|7412_  = \new_Sorter100|7312_  & \new_Sorter100|7313_ ;
  assign \new_Sorter100|7413_  = \new_Sorter100|7312_  | \new_Sorter100|7313_ ;
  assign \new_Sorter100|7414_  = \new_Sorter100|7314_  & \new_Sorter100|7315_ ;
  assign \new_Sorter100|7415_  = \new_Sorter100|7314_  | \new_Sorter100|7315_ ;
  assign \new_Sorter100|7416_  = \new_Sorter100|7316_  & \new_Sorter100|7317_ ;
  assign \new_Sorter100|7417_  = \new_Sorter100|7316_  | \new_Sorter100|7317_ ;
  assign \new_Sorter100|7418_  = \new_Sorter100|7318_  & \new_Sorter100|7319_ ;
  assign \new_Sorter100|7419_  = \new_Sorter100|7318_  | \new_Sorter100|7319_ ;
  assign \new_Sorter100|7420_  = \new_Sorter100|7320_  & \new_Sorter100|7321_ ;
  assign \new_Sorter100|7421_  = \new_Sorter100|7320_  | \new_Sorter100|7321_ ;
  assign \new_Sorter100|7422_  = \new_Sorter100|7322_  & \new_Sorter100|7323_ ;
  assign \new_Sorter100|7423_  = \new_Sorter100|7322_  | \new_Sorter100|7323_ ;
  assign \new_Sorter100|7424_  = \new_Sorter100|7324_  & \new_Sorter100|7325_ ;
  assign \new_Sorter100|7425_  = \new_Sorter100|7324_  | \new_Sorter100|7325_ ;
  assign \new_Sorter100|7426_  = \new_Sorter100|7326_  & \new_Sorter100|7327_ ;
  assign \new_Sorter100|7427_  = \new_Sorter100|7326_  | \new_Sorter100|7327_ ;
  assign \new_Sorter100|7428_  = \new_Sorter100|7328_  & \new_Sorter100|7329_ ;
  assign \new_Sorter100|7429_  = \new_Sorter100|7328_  | \new_Sorter100|7329_ ;
  assign \new_Sorter100|7430_  = \new_Sorter100|7330_  & \new_Sorter100|7331_ ;
  assign \new_Sorter100|7431_  = \new_Sorter100|7330_  | \new_Sorter100|7331_ ;
  assign \new_Sorter100|7432_  = \new_Sorter100|7332_  & \new_Sorter100|7333_ ;
  assign \new_Sorter100|7433_  = \new_Sorter100|7332_  | \new_Sorter100|7333_ ;
  assign \new_Sorter100|7434_  = \new_Sorter100|7334_  & \new_Sorter100|7335_ ;
  assign \new_Sorter100|7435_  = \new_Sorter100|7334_  | \new_Sorter100|7335_ ;
  assign \new_Sorter100|7436_  = \new_Sorter100|7336_  & \new_Sorter100|7337_ ;
  assign \new_Sorter100|7437_  = \new_Sorter100|7336_  | \new_Sorter100|7337_ ;
  assign \new_Sorter100|7438_  = \new_Sorter100|7338_  & \new_Sorter100|7339_ ;
  assign \new_Sorter100|7439_  = \new_Sorter100|7338_  | \new_Sorter100|7339_ ;
  assign \new_Sorter100|7440_  = \new_Sorter100|7340_  & \new_Sorter100|7341_ ;
  assign \new_Sorter100|7441_  = \new_Sorter100|7340_  | \new_Sorter100|7341_ ;
  assign \new_Sorter100|7442_  = \new_Sorter100|7342_  & \new_Sorter100|7343_ ;
  assign \new_Sorter100|7443_  = \new_Sorter100|7342_  | \new_Sorter100|7343_ ;
  assign \new_Sorter100|7444_  = \new_Sorter100|7344_  & \new_Sorter100|7345_ ;
  assign \new_Sorter100|7445_  = \new_Sorter100|7344_  | \new_Sorter100|7345_ ;
  assign \new_Sorter100|7446_  = \new_Sorter100|7346_  & \new_Sorter100|7347_ ;
  assign \new_Sorter100|7447_  = \new_Sorter100|7346_  | \new_Sorter100|7347_ ;
  assign \new_Sorter100|7448_  = \new_Sorter100|7348_  & \new_Sorter100|7349_ ;
  assign \new_Sorter100|7449_  = \new_Sorter100|7348_  | \new_Sorter100|7349_ ;
  assign \new_Sorter100|7450_  = \new_Sorter100|7350_  & \new_Sorter100|7351_ ;
  assign \new_Sorter100|7451_  = \new_Sorter100|7350_  | \new_Sorter100|7351_ ;
  assign \new_Sorter100|7452_  = \new_Sorter100|7352_  & \new_Sorter100|7353_ ;
  assign \new_Sorter100|7453_  = \new_Sorter100|7352_  | \new_Sorter100|7353_ ;
  assign \new_Sorter100|7454_  = \new_Sorter100|7354_  & \new_Sorter100|7355_ ;
  assign \new_Sorter100|7455_  = \new_Sorter100|7354_  | \new_Sorter100|7355_ ;
  assign \new_Sorter100|7456_  = \new_Sorter100|7356_  & \new_Sorter100|7357_ ;
  assign \new_Sorter100|7457_  = \new_Sorter100|7356_  | \new_Sorter100|7357_ ;
  assign \new_Sorter100|7458_  = \new_Sorter100|7358_  & \new_Sorter100|7359_ ;
  assign \new_Sorter100|7459_  = \new_Sorter100|7358_  | \new_Sorter100|7359_ ;
  assign \new_Sorter100|7460_  = \new_Sorter100|7360_  & \new_Sorter100|7361_ ;
  assign \new_Sorter100|7461_  = \new_Sorter100|7360_  | \new_Sorter100|7361_ ;
  assign \new_Sorter100|7462_  = \new_Sorter100|7362_  & \new_Sorter100|7363_ ;
  assign \new_Sorter100|7463_  = \new_Sorter100|7362_  | \new_Sorter100|7363_ ;
  assign \new_Sorter100|7464_  = \new_Sorter100|7364_  & \new_Sorter100|7365_ ;
  assign \new_Sorter100|7465_  = \new_Sorter100|7364_  | \new_Sorter100|7365_ ;
  assign \new_Sorter100|7466_  = \new_Sorter100|7366_  & \new_Sorter100|7367_ ;
  assign \new_Sorter100|7467_  = \new_Sorter100|7366_  | \new_Sorter100|7367_ ;
  assign \new_Sorter100|7468_  = \new_Sorter100|7368_  & \new_Sorter100|7369_ ;
  assign \new_Sorter100|7469_  = \new_Sorter100|7368_  | \new_Sorter100|7369_ ;
  assign \new_Sorter100|7470_  = \new_Sorter100|7370_  & \new_Sorter100|7371_ ;
  assign \new_Sorter100|7471_  = \new_Sorter100|7370_  | \new_Sorter100|7371_ ;
  assign \new_Sorter100|7472_  = \new_Sorter100|7372_  & \new_Sorter100|7373_ ;
  assign \new_Sorter100|7473_  = \new_Sorter100|7372_  | \new_Sorter100|7373_ ;
  assign \new_Sorter100|7474_  = \new_Sorter100|7374_  & \new_Sorter100|7375_ ;
  assign \new_Sorter100|7475_  = \new_Sorter100|7374_  | \new_Sorter100|7375_ ;
  assign \new_Sorter100|7476_  = \new_Sorter100|7376_  & \new_Sorter100|7377_ ;
  assign \new_Sorter100|7477_  = \new_Sorter100|7376_  | \new_Sorter100|7377_ ;
  assign \new_Sorter100|7478_  = \new_Sorter100|7378_  & \new_Sorter100|7379_ ;
  assign \new_Sorter100|7479_  = \new_Sorter100|7378_  | \new_Sorter100|7379_ ;
  assign \new_Sorter100|7480_  = \new_Sorter100|7380_  & \new_Sorter100|7381_ ;
  assign \new_Sorter100|7481_  = \new_Sorter100|7380_  | \new_Sorter100|7381_ ;
  assign \new_Sorter100|7482_  = \new_Sorter100|7382_  & \new_Sorter100|7383_ ;
  assign \new_Sorter100|7483_  = \new_Sorter100|7382_  | \new_Sorter100|7383_ ;
  assign \new_Sorter100|7484_  = \new_Sorter100|7384_  & \new_Sorter100|7385_ ;
  assign \new_Sorter100|7485_  = \new_Sorter100|7384_  | \new_Sorter100|7385_ ;
  assign \new_Sorter100|7486_  = \new_Sorter100|7386_  & \new_Sorter100|7387_ ;
  assign \new_Sorter100|7487_  = \new_Sorter100|7386_  | \new_Sorter100|7387_ ;
  assign \new_Sorter100|7488_  = \new_Sorter100|7388_  & \new_Sorter100|7389_ ;
  assign \new_Sorter100|7489_  = \new_Sorter100|7388_  | \new_Sorter100|7389_ ;
  assign \new_Sorter100|7490_  = \new_Sorter100|7390_  & \new_Sorter100|7391_ ;
  assign \new_Sorter100|7491_  = \new_Sorter100|7390_  | \new_Sorter100|7391_ ;
  assign \new_Sorter100|7492_  = \new_Sorter100|7392_  & \new_Sorter100|7393_ ;
  assign \new_Sorter100|7493_  = \new_Sorter100|7392_  | \new_Sorter100|7393_ ;
  assign \new_Sorter100|7494_  = \new_Sorter100|7394_  & \new_Sorter100|7395_ ;
  assign \new_Sorter100|7495_  = \new_Sorter100|7394_  | \new_Sorter100|7395_ ;
  assign \new_Sorter100|7496_  = \new_Sorter100|7396_  & \new_Sorter100|7397_ ;
  assign \new_Sorter100|7497_  = \new_Sorter100|7396_  | \new_Sorter100|7397_ ;
  assign \new_Sorter100|7498_  = \new_Sorter100|7398_  & \new_Sorter100|7399_ ;
  assign \new_Sorter100|7499_  = \new_Sorter100|7398_  | \new_Sorter100|7399_ ;
  assign \new_Sorter100|7500_  = \new_Sorter100|7400_ ;
  assign \new_Sorter100|7599_  = \new_Sorter100|7499_ ;
  assign \new_Sorter100|7501_  = \new_Sorter100|7401_  & \new_Sorter100|7402_ ;
  assign \new_Sorter100|7502_  = \new_Sorter100|7401_  | \new_Sorter100|7402_ ;
  assign \new_Sorter100|7503_  = \new_Sorter100|7403_  & \new_Sorter100|7404_ ;
  assign \new_Sorter100|7504_  = \new_Sorter100|7403_  | \new_Sorter100|7404_ ;
  assign \new_Sorter100|7505_  = \new_Sorter100|7405_  & \new_Sorter100|7406_ ;
  assign \new_Sorter100|7506_  = \new_Sorter100|7405_  | \new_Sorter100|7406_ ;
  assign \new_Sorter100|7507_  = \new_Sorter100|7407_  & \new_Sorter100|7408_ ;
  assign \new_Sorter100|7508_  = \new_Sorter100|7407_  | \new_Sorter100|7408_ ;
  assign \new_Sorter100|7509_  = \new_Sorter100|7409_  & \new_Sorter100|7410_ ;
  assign \new_Sorter100|7510_  = \new_Sorter100|7409_  | \new_Sorter100|7410_ ;
  assign \new_Sorter100|7511_  = \new_Sorter100|7411_  & \new_Sorter100|7412_ ;
  assign \new_Sorter100|7512_  = \new_Sorter100|7411_  | \new_Sorter100|7412_ ;
  assign \new_Sorter100|7513_  = \new_Sorter100|7413_  & \new_Sorter100|7414_ ;
  assign \new_Sorter100|7514_  = \new_Sorter100|7413_  | \new_Sorter100|7414_ ;
  assign \new_Sorter100|7515_  = \new_Sorter100|7415_  & \new_Sorter100|7416_ ;
  assign \new_Sorter100|7516_  = \new_Sorter100|7415_  | \new_Sorter100|7416_ ;
  assign \new_Sorter100|7517_  = \new_Sorter100|7417_  & \new_Sorter100|7418_ ;
  assign \new_Sorter100|7518_  = \new_Sorter100|7417_  | \new_Sorter100|7418_ ;
  assign \new_Sorter100|7519_  = \new_Sorter100|7419_  & \new_Sorter100|7420_ ;
  assign \new_Sorter100|7520_  = \new_Sorter100|7419_  | \new_Sorter100|7420_ ;
  assign \new_Sorter100|7521_  = \new_Sorter100|7421_  & \new_Sorter100|7422_ ;
  assign \new_Sorter100|7522_  = \new_Sorter100|7421_  | \new_Sorter100|7422_ ;
  assign \new_Sorter100|7523_  = \new_Sorter100|7423_  & \new_Sorter100|7424_ ;
  assign \new_Sorter100|7524_  = \new_Sorter100|7423_  | \new_Sorter100|7424_ ;
  assign \new_Sorter100|7525_  = \new_Sorter100|7425_  & \new_Sorter100|7426_ ;
  assign \new_Sorter100|7526_  = \new_Sorter100|7425_  | \new_Sorter100|7426_ ;
  assign \new_Sorter100|7527_  = \new_Sorter100|7427_  & \new_Sorter100|7428_ ;
  assign \new_Sorter100|7528_  = \new_Sorter100|7427_  | \new_Sorter100|7428_ ;
  assign \new_Sorter100|7529_  = \new_Sorter100|7429_  & \new_Sorter100|7430_ ;
  assign \new_Sorter100|7530_  = \new_Sorter100|7429_  | \new_Sorter100|7430_ ;
  assign \new_Sorter100|7531_  = \new_Sorter100|7431_  & \new_Sorter100|7432_ ;
  assign \new_Sorter100|7532_  = \new_Sorter100|7431_  | \new_Sorter100|7432_ ;
  assign \new_Sorter100|7533_  = \new_Sorter100|7433_  & \new_Sorter100|7434_ ;
  assign \new_Sorter100|7534_  = \new_Sorter100|7433_  | \new_Sorter100|7434_ ;
  assign \new_Sorter100|7535_  = \new_Sorter100|7435_  & \new_Sorter100|7436_ ;
  assign \new_Sorter100|7536_  = \new_Sorter100|7435_  | \new_Sorter100|7436_ ;
  assign \new_Sorter100|7537_  = \new_Sorter100|7437_  & \new_Sorter100|7438_ ;
  assign \new_Sorter100|7538_  = \new_Sorter100|7437_  | \new_Sorter100|7438_ ;
  assign \new_Sorter100|7539_  = \new_Sorter100|7439_  & \new_Sorter100|7440_ ;
  assign \new_Sorter100|7540_  = \new_Sorter100|7439_  | \new_Sorter100|7440_ ;
  assign \new_Sorter100|7541_  = \new_Sorter100|7441_  & \new_Sorter100|7442_ ;
  assign \new_Sorter100|7542_  = \new_Sorter100|7441_  | \new_Sorter100|7442_ ;
  assign \new_Sorter100|7543_  = \new_Sorter100|7443_  & \new_Sorter100|7444_ ;
  assign \new_Sorter100|7544_  = \new_Sorter100|7443_  | \new_Sorter100|7444_ ;
  assign \new_Sorter100|7545_  = \new_Sorter100|7445_  & \new_Sorter100|7446_ ;
  assign \new_Sorter100|7546_  = \new_Sorter100|7445_  | \new_Sorter100|7446_ ;
  assign \new_Sorter100|7547_  = \new_Sorter100|7447_  & \new_Sorter100|7448_ ;
  assign \new_Sorter100|7548_  = \new_Sorter100|7447_  | \new_Sorter100|7448_ ;
  assign \new_Sorter100|7549_  = \new_Sorter100|7449_  & \new_Sorter100|7450_ ;
  assign \new_Sorter100|7550_  = \new_Sorter100|7449_  | \new_Sorter100|7450_ ;
  assign \new_Sorter100|7551_  = \new_Sorter100|7451_  & \new_Sorter100|7452_ ;
  assign \new_Sorter100|7552_  = \new_Sorter100|7451_  | \new_Sorter100|7452_ ;
  assign \new_Sorter100|7553_  = \new_Sorter100|7453_  & \new_Sorter100|7454_ ;
  assign \new_Sorter100|7554_  = \new_Sorter100|7453_  | \new_Sorter100|7454_ ;
  assign \new_Sorter100|7555_  = \new_Sorter100|7455_  & \new_Sorter100|7456_ ;
  assign \new_Sorter100|7556_  = \new_Sorter100|7455_  | \new_Sorter100|7456_ ;
  assign \new_Sorter100|7557_  = \new_Sorter100|7457_  & \new_Sorter100|7458_ ;
  assign \new_Sorter100|7558_  = \new_Sorter100|7457_  | \new_Sorter100|7458_ ;
  assign \new_Sorter100|7559_  = \new_Sorter100|7459_  & \new_Sorter100|7460_ ;
  assign \new_Sorter100|7560_  = \new_Sorter100|7459_  | \new_Sorter100|7460_ ;
  assign \new_Sorter100|7561_  = \new_Sorter100|7461_  & \new_Sorter100|7462_ ;
  assign \new_Sorter100|7562_  = \new_Sorter100|7461_  | \new_Sorter100|7462_ ;
  assign \new_Sorter100|7563_  = \new_Sorter100|7463_  & \new_Sorter100|7464_ ;
  assign \new_Sorter100|7564_  = \new_Sorter100|7463_  | \new_Sorter100|7464_ ;
  assign \new_Sorter100|7565_  = \new_Sorter100|7465_  & \new_Sorter100|7466_ ;
  assign \new_Sorter100|7566_  = \new_Sorter100|7465_  | \new_Sorter100|7466_ ;
  assign \new_Sorter100|7567_  = \new_Sorter100|7467_  & \new_Sorter100|7468_ ;
  assign \new_Sorter100|7568_  = \new_Sorter100|7467_  | \new_Sorter100|7468_ ;
  assign \new_Sorter100|7569_  = \new_Sorter100|7469_  & \new_Sorter100|7470_ ;
  assign \new_Sorter100|7570_  = \new_Sorter100|7469_  | \new_Sorter100|7470_ ;
  assign \new_Sorter100|7571_  = \new_Sorter100|7471_  & \new_Sorter100|7472_ ;
  assign \new_Sorter100|7572_  = \new_Sorter100|7471_  | \new_Sorter100|7472_ ;
  assign \new_Sorter100|7573_  = \new_Sorter100|7473_  & \new_Sorter100|7474_ ;
  assign \new_Sorter100|7574_  = \new_Sorter100|7473_  | \new_Sorter100|7474_ ;
  assign \new_Sorter100|7575_  = \new_Sorter100|7475_  & \new_Sorter100|7476_ ;
  assign \new_Sorter100|7576_  = \new_Sorter100|7475_  | \new_Sorter100|7476_ ;
  assign \new_Sorter100|7577_  = \new_Sorter100|7477_  & \new_Sorter100|7478_ ;
  assign \new_Sorter100|7578_  = \new_Sorter100|7477_  | \new_Sorter100|7478_ ;
  assign \new_Sorter100|7579_  = \new_Sorter100|7479_  & \new_Sorter100|7480_ ;
  assign \new_Sorter100|7580_  = \new_Sorter100|7479_  | \new_Sorter100|7480_ ;
  assign \new_Sorter100|7581_  = \new_Sorter100|7481_  & \new_Sorter100|7482_ ;
  assign \new_Sorter100|7582_  = \new_Sorter100|7481_  | \new_Sorter100|7482_ ;
  assign \new_Sorter100|7583_  = \new_Sorter100|7483_  & \new_Sorter100|7484_ ;
  assign \new_Sorter100|7584_  = \new_Sorter100|7483_  | \new_Sorter100|7484_ ;
  assign \new_Sorter100|7585_  = \new_Sorter100|7485_  & \new_Sorter100|7486_ ;
  assign \new_Sorter100|7586_  = \new_Sorter100|7485_  | \new_Sorter100|7486_ ;
  assign \new_Sorter100|7587_  = \new_Sorter100|7487_  & \new_Sorter100|7488_ ;
  assign \new_Sorter100|7588_  = \new_Sorter100|7487_  | \new_Sorter100|7488_ ;
  assign \new_Sorter100|7589_  = \new_Sorter100|7489_  & \new_Sorter100|7490_ ;
  assign \new_Sorter100|7590_  = \new_Sorter100|7489_  | \new_Sorter100|7490_ ;
  assign \new_Sorter100|7591_  = \new_Sorter100|7491_  & \new_Sorter100|7492_ ;
  assign \new_Sorter100|7592_  = \new_Sorter100|7491_  | \new_Sorter100|7492_ ;
  assign \new_Sorter100|7593_  = \new_Sorter100|7493_  & \new_Sorter100|7494_ ;
  assign \new_Sorter100|7594_  = \new_Sorter100|7493_  | \new_Sorter100|7494_ ;
  assign \new_Sorter100|7595_  = \new_Sorter100|7495_  & \new_Sorter100|7496_ ;
  assign \new_Sorter100|7596_  = \new_Sorter100|7495_  | \new_Sorter100|7496_ ;
  assign \new_Sorter100|7597_  = \new_Sorter100|7497_  & \new_Sorter100|7498_ ;
  assign \new_Sorter100|7598_  = \new_Sorter100|7497_  | \new_Sorter100|7498_ ;
  assign \new_Sorter100|7600_  = \new_Sorter100|7500_  & \new_Sorter100|7501_ ;
  assign \new_Sorter100|7601_  = \new_Sorter100|7500_  | \new_Sorter100|7501_ ;
  assign \new_Sorter100|7602_  = \new_Sorter100|7502_  & \new_Sorter100|7503_ ;
  assign \new_Sorter100|7603_  = \new_Sorter100|7502_  | \new_Sorter100|7503_ ;
  assign \new_Sorter100|7604_  = \new_Sorter100|7504_  & \new_Sorter100|7505_ ;
  assign \new_Sorter100|7605_  = \new_Sorter100|7504_  | \new_Sorter100|7505_ ;
  assign \new_Sorter100|7606_  = \new_Sorter100|7506_  & \new_Sorter100|7507_ ;
  assign \new_Sorter100|7607_  = \new_Sorter100|7506_  | \new_Sorter100|7507_ ;
  assign \new_Sorter100|7608_  = \new_Sorter100|7508_  & \new_Sorter100|7509_ ;
  assign \new_Sorter100|7609_  = \new_Sorter100|7508_  | \new_Sorter100|7509_ ;
  assign \new_Sorter100|7610_  = \new_Sorter100|7510_  & \new_Sorter100|7511_ ;
  assign \new_Sorter100|7611_  = \new_Sorter100|7510_  | \new_Sorter100|7511_ ;
  assign \new_Sorter100|7612_  = \new_Sorter100|7512_  & \new_Sorter100|7513_ ;
  assign \new_Sorter100|7613_  = \new_Sorter100|7512_  | \new_Sorter100|7513_ ;
  assign \new_Sorter100|7614_  = \new_Sorter100|7514_  & \new_Sorter100|7515_ ;
  assign \new_Sorter100|7615_  = \new_Sorter100|7514_  | \new_Sorter100|7515_ ;
  assign \new_Sorter100|7616_  = \new_Sorter100|7516_  & \new_Sorter100|7517_ ;
  assign \new_Sorter100|7617_  = \new_Sorter100|7516_  | \new_Sorter100|7517_ ;
  assign \new_Sorter100|7618_  = \new_Sorter100|7518_  & \new_Sorter100|7519_ ;
  assign \new_Sorter100|7619_  = \new_Sorter100|7518_  | \new_Sorter100|7519_ ;
  assign \new_Sorter100|7620_  = \new_Sorter100|7520_  & \new_Sorter100|7521_ ;
  assign \new_Sorter100|7621_  = \new_Sorter100|7520_  | \new_Sorter100|7521_ ;
  assign \new_Sorter100|7622_  = \new_Sorter100|7522_  & \new_Sorter100|7523_ ;
  assign \new_Sorter100|7623_  = \new_Sorter100|7522_  | \new_Sorter100|7523_ ;
  assign \new_Sorter100|7624_  = \new_Sorter100|7524_  & \new_Sorter100|7525_ ;
  assign \new_Sorter100|7625_  = \new_Sorter100|7524_  | \new_Sorter100|7525_ ;
  assign \new_Sorter100|7626_  = \new_Sorter100|7526_  & \new_Sorter100|7527_ ;
  assign \new_Sorter100|7627_  = \new_Sorter100|7526_  | \new_Sorter100|7527_ ;
  assign \new_Sorter100|7628_  = \new_Sorter100|7528_  & \new_Sorter100|7529_ ;
  assign \new_Sorter100|7629_  = \new_Sorter100|7528_  | \new_Sorter100|7529_ ;
  assign \new_Sorter100|7630_  = \new_Sorter100|7530_  & \new_Sorter100|7531_ ;
  assign \new_Sorter100|7631_  = \new_Sorter100|7530_  | \new_Sorter100|7531_ ;
  assign \new_Sorter100|7632_  = \new_Sorter100|7532_  & \new_Sorter100|7533_ ;
  assign \new_Sorter100|7633_  = \new_Sorter100|7532_  | \new_Sorter100|7533_ ;
  assign \new_Sorter100|7634_  = \new_Sorter100|7534_  & \new_Sorter100|7535_ ;
  assign \new_Sorter100|7635_  = \new_Sorter100|7534_  | \new_Sorter100|7535_ ;
  assign \new_Sorter100|7636_  = \new_Sorter100|7536_  & \new_Sorter100|7537_ ;
  assign \new_Sorter100|7637_  = \new_Sorter100|7536_  | \new_Sorter100|7537_ ;
  assign \new_Sorter100|7638_  = \new_Sorter100|7538_  & \new_Sorter100|7539_ ;
  assign \new_Sorter100|7639_  = \new_Sorter100|7538_  | \new_Sorter100|7539_ ;
  assign \new_Sorter100|7640_  = \new_Sorter100|7540_  & \new_Sorter100|7541_ ;
  assign \new_Sorter100|7641_  = \new_Sorter100|7540_  | \new_Sorter100|7541_ ;
  assign \new_Sorter100|7642_  = \new_Sorter100|7542_  & \new_Sorter100|7543_ ;
  assign \new_Sorter100|7643_  = \new_Sorter100|7542_  | \new_Sorter100|7543_ ;
  assign \new_Sorter100|7644_  = \new_Sorter100|7544_  & \new_Sorter100|7545_ ;
  assign \new_Sorter100|7645_  = \new_Sorter100|7544_  | \new_Sorter100|7545_ ;
  assign \new_Sorter100|7646_  = \new_Sorter100|7546_  & \new_Sorter100|7547_ ;
  assign \new_Sorter100|7647_  = \new_Sorter100|7546_  | \new_Sorter100|7547_ ;
  assign \new_Sorter100|7648_  = \new_Sorter100|7548_  & \new_Sorter100|7549_ ;
  assign \new_Sorter100|7649_  = \new_Sorter100|7548_  | \new_Sorter100|7549_ ;
  assign \new_Sorter100|7650_  = \new_Sorter100|7550_  & \new_Sorter100|7551_ ;
  assign \new_Sorter100|7651_  = \new_Sorter100|7550_  | \new_Sorter100|7551_ ;
  assign \new_Sorter100|7652_  = \new_Sorter100|7552_  & \new_Sorter100|7553_ ;
  assign \new_Sorter100|7653_  = \new_Sorter100|7552_  | \new_Sorter100|7553_ ;
  assign \new_Sorter100|7654_  = \new_Sorter100|7554_  & \new_Sorter100|7555_ ;
  assign \new_Sorter100|7655_  = \new_Sorter100|7554_  | \new_Sorter100|7555_ ;
  assign \new_Sorter100|7656_  = \new_Sorter100|7556_  & \new_Sorter100|7557_ ;
  assign \new_Sorter100|7657_  = \new_Sorter100|7556_  | \new_Sorter100|7557_ ;
  assign \new_Sorter100|7658_  = \new_Sorter100|7558_  & \new_Sorter100|7559_ ;
  assign \new_Sorter100|7659_  = \new_Sorter100|7558_  | \new_Sorter100|7559_ ;
  assign \new_Sorter100|7660_  = \new_Sorter100|7560_  & \new_Sorter100|7561_ ;
  assign \new_Sorter100|7661_  = \new_Sorter100|7560_  | \new_Sorter100|7561_ ;
  assign \new_Sorter100|7662_  = \new_Sorter100|7562_  & \new_Sorter100|7563_ ;
  assign \new_Sorter100|7663_  = \new_Sorter100|7562_  | \new_Sorter100|7563_ ;
  assign \new_Sorter100|7664_  = \new_Sorter100|7564_  & \new_Sorter100|7565_ ;
  assign \new_Sorter100|7665_  = \new_Sorter100|7564_  | \new_Sorter100|7565_ ;
  assign \new_Sorter100|7666_  = \new_Sorter100|7566_  & \new_Sorter100|7567_ ;
  assign \new_Sorter100|7667_  = \new_Sorter100|7566_  | \new_Sorter100|7567_ ;
  assign \new_Sorter100|7668_  = \new_Sorter100|7568_  & \new_Sorter100|7569_ ;
  assign \new_Sorter100|7669_  = \new_Sorter100|7568_  | \new_Sorter100|7569_ ;
  assign \new_Sorter100|7670_  = \new_Sorter100|7570_  & \new_Sorter100|7571_ ;
  assign \new_Sorter100|7671_  = \new_Sorter100|7570_  | \new_Sorter100|7571_ ;
  assign \new_Sorter100|7672_  = \new_Sorter100|7572_  & \new_Sorter100|7573_ ;
  assign \new_Sorter100|7673_  = \new_Sorter100|7572_  | \new_Sorter100|7573_ ;
  assign \new_Sorter100|7674_  = \new_Sorter100|7574_  & \new_Sorter100|7575_ ;
  assign \new_Sorter100|7675_  = \new_Sorter100|7574_  | \new_Sorter100|7575_ ;
  assign \new_Sorter100|7676_  = \new_Sorter100|7576_  & \new_Sorter100|7577_ ;
  assign \new_Sorter100|7677_  = \new_Sorter100|7576_  | \new_Sorter100|7577_ ;
  assign \new_Sorter100|7678_  = \new_Sorter100|7578_  & \new_Sorter100|7579_ ;
  assign \new_Sorter100|7679_  = \new_Sorter100|7578_  | \new_Sorter100|7579_ ;
  assign \new_Sorter100|7680_  = \new_Sorter100|7580_  & \new_Sorter100|7581_ ;
  assign \new_Sorter100|7681_  = \new_Sorter100|7580_  | \new_Sorter100|7581_ ;
  assign \new_Sorter100|7682_  = \new_Sorter100|7582_  & \new_Sorter100|7583_ ;
  assign \new_Sorter100|7683_  = \new_Sorter100|7582_  | \new_Sorter100|7583_ ;
  assign \new_Sorter100|7684_  = \new_Sorter100|7584_  & \new_Sorter100|7585_ ;
  assign \new_Sorter100|7685_  = \new_Sorter100|7584_  | \new_Sorter100|7585_ ;
  assign \new_Sorter100|7686_  = \new_Sorter100|7586_  & \new_Sorter100|7587_ ;
  assign \new_Sorter100|7687_  = \new_Sorter100|7586_  | \new_Sorter100|7587_ ;
  assign \new_Sorter100|7688_  = \new_Sorter100|7588_  & \new_Sorter100|7589_ ;
  assign \new_Sorter100|7689_  = \new_Sorter100|7588_  | \new_Sorter100|7589_ ;
  assign \new_Sorter100|7690_  = \new_Sorter100|7590_  & \new_Sorter100|7591_ ;
  assign \new_Sorter100|7691_  = \new_Sorter100|7590_  | \new_Sorter100|7591_ ;
  assign \new_Sorter100|7692_  = \new_Sorter100|7592_  & \new_Sorter100|7593_ ;
  assign \new_Sorter100|7693_  = \new_Sorter100|7592_  | \new_Sorter100|7593_ ;
  assign \new_Sorter100|7694_  = \new_Sorter100|7594_  & \new_Sorter100|7595_ ;
  assign \new_Sorter100|7695_  = \new_Sorter100|7594_  | \new_Sorter100|7595_ ;
  assign \new_Sorter100|7696_  = \new_Sorter100|7596_  & \new_Sorter100|7597_ ;
  assign \new_Sorter100|7697_  = \new_Sorter100|7596_  | \new_Sorter100|7597_ ;
  assign \new_Sorter100|7698_  = \new_Sorter100|7598_  & \new_Sorter100|7599_ ;
  assign \new_Sorter100|7699_  = \new_Sorter100|7598_  | \new_Sorter100|7599_ ;
  assign \new_Sorter100|7700_  = \new_Sorter100|7600_ ;
  assign \new_Sorter100|7799_  = \new_Sorter100|7699_ ;
  assign \new_Sorter100|7701_  = \new_Sorter100|7601_  & \new_Sorter100|7602_ ;
  assign \new_Sorter100|7702_  = \new_Sorter100|7601_  | \new_Sorter100|7602_ ;
  assign \new_Sorter100|7703_  = \new_Sorter100|7603_  & \new_Sorter100|7604_ ;
  assign \new_Sorter100|7704_  = \new_Sorter100|7603_  | \new_Sorter100|7604_ ;
  assign \new_Sorter100|7705_  = \new_Sorter100|7605_  & \new_Sorter100|7606_ ;
  assign \new_Sorter100|7706_  = \new_Sorter100|7605_  | \new_Sorter100|7606_ ;
  assign \new_Sorter100|7707_  = \new_Sorter100|7607_  & \new_Sorter100|7608_ ;
  assign \new_Sorter100|7708_  = \new_Sorter100|7607_  | \new_Sorter100|7608_ ;
  assign \new_Sorter100|7709_  = \new_Sorter100|7609_  & \new_Sorter100|7610_ ;
  assign \new_Sorter100|7710_  = \new_Sorter100|7609_  | \new_Sorter100|7610_ ;
  assign \new_Sorter100|7711_  = \new_Sorter100|7611_  & \new_Sorter100|7612_ ;
  assign \new_Sorter100|7712_  = \new_Sorter100|7611_  | \new_Sorter100|7612_ ;
  assign \new_Sorter100|7713_  = \new_Sorter100|7613_  & \new_Sorter100|7614_ ;
  assign \new_Sorter100|7714_  = \new_Sorter100|7613_  | \new_Sorter100|7614_ ;
  assign \new_Sorter100|7715_  = \new_Sorter100|7615_  & \new_Sorter100|7616_ ;
  assign \new_Sorter100|7716_  = \new_Sorter100|7615_  | \new_Sorter100|7616_ ;
  assign \new_Sorter100|7717_  = \new_Sorter100|7617_  & \new_Sorter100|7618_ ;
  assign \new_Sorter100|7718_  = \new_Sorter100|7617_  | \new_Sorter100|7618_ ;
  assign \new_Sorter100|7719_  = \new_Sorter100|7619_  & \new_Sorter100|7620_ ;
  assign \new_Sorter100|7720_  = \new_Sorter100|7619_  | \new_Sorter100|7620_ ;
  assign \new_Sorter100|7721_  = \new_Sorter100|7621_  & \new_Sorter100|7622_ ;
  assign \new_Sorter100|7722_  = \new_Sorter100|7621_  | \new_Sorter100|7622_ ;
  assign \new_Sorter100|7723_  = \new_Sorter100|7623_  & \new_Sorter100|7624_ ;
  assign \new_Sorter100|7724_  = \new_Sorter100|7623_  | \new_Sorter100|7624_ ;
  assign \new_Sorter100|7725_  = \new_Sorter100|7625_  & \new_Sorter100|7626_ ;
  assign \new_Sorter100|7726_  = \new_Sorter100|7625_  | \new_Sorter100|7626_ ;
  assign \new_Sorter100|7727_  = \new_Sorter100|7627_  & \new_Sorter100|7628_ ;
  assign \new_Sorter100|7728_  = \new_Sorter100|7627_  | \new_Sorter100|7628_ ;
  assign \new_Sorter100|7729_  = \new_Sorter100|7629_  & \new_Sorter100|7630_ ;
  assign \new_Sorter100|7730_  = \new_Sorter100|7629_  | \new_Sorter100|7630_ ;
  assign \new_Sorter100|7731_  = \new_Sorter100|7631_  & \new_Sorter100|7632_ ;
  assign \new_Sorter100|7732_  = \new_Sorter100|7631_  | \new_Sorter100|7632_ ;
  assign \new_Sorter100|7733_  = \new_Sorter100|7633_  & \new_Sorter100|7634_ ;
  assign \new_Sorter100|7734_  = \new_Sorter100|7633_  | \new_Sorter100|7634_ ;
  assign \new_Sorter100|7735_  = \new_Sorter100|7635_  & \new_Sorter100|7636_ ;
  assign \new_Sorter100|7736_  = \new_Sorter100|7635_  | \new_Sorter100|7636_ ;
  assign \new_Sorter100|7737_  = \new_Sorter100|7637_  & \new_Sorter100|7638_ ;
  assign \new_Sorter100|7738_  = \new_Sorter100|7637_  | \new_Sorter100|7638_ ;
  assign \new_Sorter100|7739_  = \new_Sorter100|7639_  & \new_Sorter100|7640_ ;
  assign \new_Sorter100|7740_  = \new_Sorter100|7639_  | \new_Sorter100|7640_ ;
  assign \new_Sorter100|7741_  = \new_Sorter100|7641_  & \new_Sorter100|7642_ ;
  assign \new_Sorter100|7742_  = \new_Sorter100|7641_  | \new_Sorter100|7642_ ;
  assign \new_Sorter100|7743_  = \new_Sorter100|7643_  & \new_Sorter100|7644_ ;
  assign \new_Sorter100|7744_  = \new_Sorter100|7643_  | \new_Sorter100|7644_ ;
  assign \new_Sorter100|7745_  = \new_Sorter100|7645_  & \new_Sorter100|7646_ ;
  assign \new_Sorter100|7746_  = \new_Sorter100|7645_  | \new_Sorter100|7646_ ;
  assign \new_Sorter100|7747_  = \new_Sorter100|7647_  & \new_Sorter100|7648_ ;
  assign \new_Sorter100|7748_  = \new_Sorter100|7647_  | \new_Sorter100|7648_ ;
  assign \new_Sorter100|7749_  = \new_Sorter100|7649_  & \new_Sorter100|7650_ ;
  assign \new_Sorter100|7750_  = \new_Sorter100|7649_  | \new_Sorter100|7650_ ;
  assign \new_Sorter100|7751_  = \new_Sorter100|7651_  & \new_Sorter100|7652_ ;
  assign \new_Sorter100|7752_  = \new_Sorter100|7651_  | \new_Sorter100|7652_ ;
  assign \new_Sorter100|7753_  = \new_Sorter100|7653_  & \new_Sorter100|7654_ ;
  assign \new_Sorter100|7754_  = \new_Sorter100|7653_  | \new_Sorter100|7654_ ;
  assign \new_Sorter100|7755_  = \new_Sorter100|7655_  & \new_Sorter100|7656_ ;
  assign \new_Sorter100|7756_  = \new_Sorter100|7655_  | \new_Sorter100|7656_ ;
  assign \new_Sorter100|7757_  = \new_Sorter100|7657_  & \new_Sorter100|7658_ ;
  assign \new_Sorter100|7758_  = \new_Sorter100|7657_  | \new_Sorter100|7658_ ;
  assign \new_Sorter100|7759_  = \new_Sorter100|7659_  & \new_Sorter100|7660_ ;
  assign \new_Sorter100|7760_  = \new_Sorter100|7659_  | \new_Sorter100|7660_ ;
  assign \new_Sorter100|7761_  = \new_Sorter100|7661_  & \new_Sorter100|7662_ ;
  assign \new_Sorter100|7762_  = \new_Sorter100|7661_  | \new_Sorter100|7662_ ;
  assign \new_Sorter100|7763_  = \new_Sorter100|7663_  & \new_Sorter100|7664_ ;
  assign \new_Sorter100|7764_  = \new_Sorter100|7663_  | \new_Sorter100|7664_ ;
  assign \new_Sorter100|7765_  = \new_Sorter100|7665_  & \new_Sorter100|7666_ ;
  assign \new_Sorter100|7766_  = \new_Sorter100|7665_  | \new_Sorter100|7666_ ;
  assign \new_Sorter100|7767_  = \new_Sorter100|7667_  & \new_Sorter100|7668_ ;
  assign \new_Sorter100|7768_  = \new_Sorter100|7667_  | \new_Sorter100|7668_ ;
  assign \new_Sorter100|7769_  = \new_Sorter100|7669_  & \new_Sorter100|7670_ ;
  assign \new_Sorter100|7770_  = \new_Sorter100|7669_  | \new_Sorter100|7670_ ;
  assign \new_Sorter100|7771_  = \new_Sorter100|7671_  & \new_Sorter100|7672_ ;
  assign \new_Sorter100|7772_  = \new_Sorter100|7671_  | \new_Sorter100|7672_ ;
  assign \new_Sorter100|7773_  = \new_Sorter100|7673_  & \new_Sorter100|7674_ ;
  assign \new_Sorter100|7774_  = \new_Sorter100|7673_  | \new_Sorter100|7674_ ;
  assign \new_Sorter100|7775_  = \new_Sorter100|7675_  & \new_Sorter100|7676_ ;
  assign \new_Sorter100|7776_  = \new_Sorter100|7675_  | \new_Sorter100|7676_ ;
  assign \new_Sorter100|7777_  = \new_Sorter100|7677_  & \new_Sorter100|7678_ ;
  assign \new_Sorter100|7778_  = \new_Sorter100|7677_  | \new_Sorter100|7678_ ;
  assign \new_Sorter100|7779_  = \new_Sorter100|7679_  & \new_Sorter100|7680_ ;
  assign \new_Sorter100|7780_  = \new_Sorter100|7679_  | \new_Sorter100|7680_ ;
  assign \new_Sorter100|7781_  = \new_Sorter100|7681_  & \new_Sorter100|7682_ ;
  assign \new_Sorter100|7782_  = \new_Sorter100|7681_  | \new_Sorter100|7682_ ;
  assign \new_Sorter100|7783_  = \new_Sorter100|7683_  & \new_Sorter100|7684_ ;
  assign \new_Sorter100|7784_  = \new_Sorter100|7683_  | \new_Sorter100|7684_ ;
  assign \new_Sorter100|7785_  = \new_Sorter100|7685_  & \new_Sorter100|7686_ ;
  assign \new_Sorter100|7786_  = \new_Sorter100|7685_  | \new_Sorter100|7686_ ;
  assign \new_Sorter100|7787_  = \new_Sorter100|7687_  & \new_Sorter100|7688_ ;
  assign \new_Sorter100|7788_  = \new_Sorter100|7687_  | \new_Sorter100|7688_ ;
  assign \new_Sorter100|7789_  = \new_Sorter100|7689_  & \new_Sorter100|7690_ ;
  assign \new_Sorter100|7790_  = \new_Sorter100|7689_  | \new_Sorter100|7690_ ;
  assign \new_Sorter100|7791_  = \new_Sorter100|7691_  & \new_Sorter100|7692_ ;
  assign \new_Sorter100|7792_  = \new_Sorter100|7691_  | \new_Sorter100|7692_ ;
  assign \new_Sorter100|7793_  = \new_Sorter100|7693_  & \new_Sorter100|7694_ ;
  assign \new_Sorter100|7794_  = \new_Sorter100|7693_  | \new_Sorter100|7694_ ;
  assign \new_Sorter100|7795_  = \new_Sorter100|7695_  & \new_Sorter100|7696_ ;
  assign \new_Sorter100|7796_  = \new_Sorter100|7695_  | \new_Sorter100|7696_ ;
  assign \new_Sorter100|7797_  = \new_Sorter100|7697_  & \new_Sorter100|7698_ ;
  assign \new_Sorter100|7798_  = \new_Sorter100|7697_  | \new_Sorter100|7698_ ;
  assign \new_Sorter100|7800_  = \new_Sorter100|7700_  & \new_Sorter100|7701_ ;
  assign \new_Sorter100|7801_  = \new_Sorter100|7700_  | \new_Sorter100|7701_ ;
  assign \new_Sorter100|7802_  = \new_Sorter100|7702_  & \new_Sorter100|7703_ ;
  assign \new_Sorter100|7803_  = \new_Sorter100|7702_  | \new_Sorter100|7703_ ;
  assign \new_Sorter100|7804_  = \new_Sorter100|7704_  & \new_Sorter100|7705_ ;
  assign \new_Sorter100|7805_  = \new_Sorter100|7704_  | \new_Sorter100|7705_ ;
  assign \new_Sorter100|7806_  = \new_Sorter100|7706_  & \new_Sorter100|7707_ ;
  assign \new_Sorter100|7807_  = \new_Sorter100|7706_  | \new_Sorter100|7707_ ;
  assign \new_Sorter100|7808_  = \new_Sorter100|7708_  & \new_Sorter100|7709_ ;
  assign \new_Sorter100|7809_  = \new_Sorter100|7708_  | \new_Sorter100|7709_ ;
  assign \new_Sorter100|7810_  = \new_Sorter100|7710_  & \new_Sorter100|7711_ ;
  assign \new_Sorter100|7811_  = \new_Sorter100|7710_  | \new_Sorter100|7711_ ;
  assign \new_Sorter100|7812_  = \new_Sorter100|7712_  & \new_Sorter100|7713_ ;
  assign \new_Sorter100|7813_  = \new_Sorter100|7712_  | \new_Sorter100|7713_ ;
  assign \new_Sorter100|7814_  = \new_Sorter100|7714_  & \new_Sorter100|7715_ ;
  assign \new_Sorter100|7815_  = \new_Sorter100|7714_  | \new_Sorter100|7715_ ;
  assign \new_Sorter100|7816_  = \new_Sorter100|7716_  & \new_Sorter100|7717_ ;
  assign \new_Sorter100|7817_  = \new_Sorter100|7716_  | \new_Sorter100|7717_ ;
  assign \new_Sorter100|7818_  = \new_Sorter100|7718_  & \new_Sorter100|7719_ ;
  assign \new_Sorter100|7819_  = \new_Sorter100|7718_  | \new_Sorter100|7719_ ;
  assign \new_Sorter100|7820_  = \new_Sorter100|7720_  & \new_Sorter100|7721_ ;
  assign \new_Sorter100|7821_  = \new_Sorter100|7720_  | \new_Sorter100|7721_ ;
  assign \new_Sorter100|7822_  = \new_Sorter100|7722_  & \new_Sorter100|7723_ ;
  assign \new_Sorter100|7823_  = \new_Sorter100|7722_  | \new_Sorter100|7723_ ;
  assign \new_Sorter100|7824_  = \new_Sorter100|7724_  & \new_Sorter100|7725_ ;
  assign \new_Sorter100|7825_  = \new_Sorter100|7724_  | \new_Sorter100|7725_ ;
  assign \new_Sorter100|7826_  = \new_Sorter100|7726_  & \new_Sorter100|7727_ ;
  assign \new_Sorter100|7827_  = \new_Sorter100|7726_  | \new_Sorter100|7727_ ;
  assign \new_Sorter100|7828_  = \new_Sorter100|7728_  & \new_Sorter100|7729_ ;
  assign \new_Sorter100|7829_  = \new_Sorter100|7728_  | \new_Sorter100|7729_ ;
  assign \new_Sorter100|7830_  = \new_Sorter100|7730_  & \new_Sorter100|7731_ ;
  assign \new_Sorter100|7831_  = \new_Sorter100|7730_  | \new_Sorter100|7731_ ;
  assign \new_Sorter100|7832_  = \new_Sorter100|7732_  & \new_Sorter100|7733_ ;
  assign \new_Sorter100|7833_  = \new_Sorter100|7732_  | \new_Sorter100|7733_ ;
  assign \new_Sorter100|7834_  = \new_Sorter100|7734_  & \new_Sorter100|7735_ ;
  assign \new_Sorter100|7835_  = \new_Sorter100|7734_  | \new_Sorter100|7735_ ;
  assign \new_Sorter100|7836_  = \new_Sorter100|7736_  & \new_Sorter100|7737_ ;
  assign \new_Sorter100|7837_  = \new_Sorter100|7736_  | \new_Sorter100|7737_ ;
  assign \new_Sorter100|7838_  = \new_Sorter100|7738_  & \new_Sorter100|7739_ ;
  assign \new_Sorter100|7839_  = \new_Sorter100|7738_  | \new_Sorter100|7739_ ;
  assign \new_Sorter100|7840_  = \new_Sorter100|7740_  & \new_Sorter100|7741_ ;
  assign \new_Sorter100|7841_  = \new_Sorter100|7740_  | \new_Sorter100|7741_ ;
  assign \new_Sorter100|7842_  = \new_Sorter100|7742_  & \new_Sorter100|7743_ ;
  assign \new_Sorter100|7843_  = \new_Sorter100|7742_  | \new_Sorter100|7743_ ;
  assign \new_Sorter100|7844_  = \new_Sorter100|7744_  & \new_Sorter100|7745_ ;
  assign \new_Sorter100|7845_  = \new_Sorter100|7744_  | \new_Sorter100|7745_ ;
  assign \new_Sorter100|7846_  = \new_Sorter100|7746_  & \new_Sorter100|7747_ ;
  assign \new_Sorter100|7847_  = \new_Sorter100|7746_  | \new_Sorter100|7747_ ;
  assign \new_Sorter100|7848_  = \new_Sorter100|7748_  & \new_Sorter100|7749_ ;
  assign \new_Sorter100|7849_  = \new_Sorter100|7748_  | \new_Sorter100|7749_ ;
  assign \new_Sorter100|7850_  = \new_Sorter100|7750_  & \new_Sorter100|7751_ ;
  assign \new_Sorter100|7851_  = \new_Sorter100|7750_  | \new_Sorter100|7751_ ;
  assign \new_Sorter100|7852_  = \new_Sorter100|7752_  & \new_Sorter100|7753_ ;
  assign \new_Sorter100|7853_  = \new_Sorter100|7752_  | \new_Sorter100|7753_ ;
  assign \new_Sorter100|7854_  = \new_Sorter100|7754_  & \new_Sorter100|7755_ ;
  assign \new_Sorter100|7855_  = \new_Sorter100|7754_  | \new_Sorter100|7755_ ;
  assign \new_Sorter100|7856_  = \new_Sorter100|7756_  & \new_Sorter100|7757_ ;
  assign \new_Sorter100|7857_  = \new_Sorter100|7756_  | \new_Sorter100|7757_ ;
  assign \new_Sorter100|7858_  = \new_Sorter100|7758_  & \new_Sorter100|7759_ ;
  assign \new_Sorter100|7859_  = \new_Sorter100|7758_  | \new_Sorter100|7759_ ;
  assign \new_Sorter100|7860_  = \new_Sorter100|7760_  & \new_Sorter100|7761_ ;
  assign \new_Sorter100|7861_  = \new_Sorter100|7760_  | \new_Sorter100|7761_ ;
  assign \new_Sorter100|7862_  = \new_Sorter100|7762_  & \new_Sorter100|7763_ ;
  assign \new_Sorter100|7863_  = \new_Sorter100|7762_  | \new_Sorter100|7763_ ;
  assign \new_Sorter100|7864_  = \new_Sorter100|7764_  & \new_Sorter100|7765_ ;
  assign \new_Sorter100|7865_  = \new_Sorter100|7764_  | \new_Sorter100|7765_ ;
  assign \new_Sorter100|7866_  = \new_Sorter100|7766_  & \new_Sorter100|7767_ ;
  assign \new_Sorter100|7867_  = \new_Sorter100|7766_  | \new_Sorter100|7767_ ;
  assign \new_Sorter100|7868_  = \new_Sorter100|7768_  & \new_Sorter100|7769_ ;
  assign \new_Sorter100|7869_  = \new_Sorter100|7768_  | \new_Sorter100|7769_ ;
  assign \new_Sorter100|7870_  = \new_Sorter100|7770_  & \new_Sorter100|7771_ ;
  assign \new_Sorter100|7871_  = \new_Sorter100|7770_  | \new_Sorter100|7771_ ;
  assign \new_Sorter100|7872_  = \new_Sorter100|7772_  & \new_Sorter100|7773_ ;
  assign \new_Sorter100|7873_  = \new_Sorter100|7772_  | \new_Sorter100|7773_ ;
  assign \new_Sorter100|7874_  = \new_Sorter100|7774_  & \new_Sorter100|7775_ ;
  assign \new_Sorter100|7875_  = \new_Sorter100|7774_  | \new_Sorter100|7775_ ;
  assign \new_Sorter100|7876_  = \new_Sorter100|7776_  & \new_Sorter100|7777_ ;
  assign \new_Sorter100|7877_  = \new_Sorter100|7776_  | \new_Sorter100|7777_ ;
  assign \new_Sorter100|7878_  = \new_Sorter100|7778_  & \new_Sorter100|7779_ ;
  assign \new_Sorter100|7879_  = \new_Sorter100|7778_  | \new_Sorter100|7779_ ;
  assign \new_Sorter100|7880_  = \new_Sorter100|7780_  & \new_Sorter100|7781_ ;
  assign \new_Sorter100|7881_  = \new_Sorter100|7780_  | \new_Sorter100|7781_ ;
  assign \new_Sorter100|7882_  = \new_Sorter100|7782_  & \new_Sorter100|7783_ ;
  assign \new_Sorter100|7883_  = \new_Sorter100|7782_  | \new_Sorter100|7783_ ;
  assign \new_Sorter100|7884_  = \new_Sorter100|7784_  & \new_Sorter100|7785_ ;
  assign \new_Sorter100|7885_  = \new_Sorter100|7784_  | \new_Sorter100|7785_ ;
  assign \new_Sorter100|7886_  = \new_Sorter100|7786_  & \new_Sorter100|7787_ ;
  assign \new_Sorter100|7887_  = \new_Sorter100|7786_  | \new_Sorter100|7787_ ;
  assign \new_Sorter100|7888_  = \new_Sorter100|7788_  & \new_Sorter100|7789_ ;
  assign \new_Sorter100|7889_  = \new_Sorter100|7788_  | \new_Sorter100|7789_ ;
  assign \new_Sorter100|7890_  = \new_Sorter100|7790_  & \new_Sorter100|7791_ ;
  assign \new_Sorter100|7891_  = \new_Sorter100|7790_  | \new_Sorter100|7791_ ;
  assign \new_Sorter100|7892_  = \new_Sorter100|7792_  & \new_Sorter100|7793_ ;
  assign \new_Sorter100|7893_  = \new_Sorter100|7792_  | \new_Sorter100|7793_ ;
  assign \new_Sorter100|7894_  = \new_Sorter100|7794_  & \new_Sorter100|7795_ ;
  assign \new_Sorter100|7895_  = \new_Sorter100|7794_  | \new_Sorter100|7795_ ;
  assign \new_Sorter100|7896_  = \new_Sorter100|7796_  & \new_Sorter100|7797_ ;
  assign \new_Sorter100|7897_  = \new_Sorter100|7796_  | \new_Sorter100|7797_ ;
  assign \new_Sorter100|7898_  = \new_Sorter100|7798_  & \new_Sorter100|7799_ ;
  assign \new_Sorter100|7899_  = \new_Sorter100|7798_  | \new_Sorter100|7799_ ;
  assign \new_Sorter100|7900_  = \new_Sorter100|7800_ ;
  assign \new_Sorter100|7999_  = \new_Sorter100|7899_ ;
  assign \new_Sorter100|7901_  = \new_Sorter100|7801_  & \new_Sorter100|7802_ ;
  assign \new_Sorter100|7902_  = \new_Sorter100|7801_  | \new_Sorter100|7802_ ;
  assign \new_Sorter100|7903_  = \new_Sorter100|7803_  & \new_Sorter100|7804_ ;
  assign \new_Sorter100|7904_  = \new_Sorter100|7803_  | \new_Sorter100|7804_ ;
  assign \new_Sorter100|7905_  = \new_Sorter100|7805_  & \new_Sorter100|7806_ ;
  assign \new_Sorter100|7906_  = \new_Sorter100|7805_  | \new_Sorter100|7806_ ;
  assign \new_Sorter100|7907_  = \new_Sorter100|7807_  & \new_Sorter100|7808_ ;
  assign \new_Sorter100|7908_  = \new_Sorter100|7807_  | \new_Sorter100|7808_ ;
  assign \new_Sorter100|7909_  = \new_Sorter100|7809_  & \new_Sorter100|7810_ ;
  assign \new_Sorter100|7910_  = \new_Sorter100|7809_  | \new_Sorter100|7810_ ;
  assign \new_Sorter100|7911_  = \new_Sorter100|7811_  & \new_Sorter100|7812_ ;
  assign \new_Sorter100|7912_  = \new_Sorter100|7811_  | \new_Sorter100|7812_ ;
  assign \new_Sorter100|7913_  = \new_Sorter100|7813_  & \new_Sorter100|7814_ ;
  assign \new_Sorter100|7914_  = \new_Sorter100|7813_  | \new_Sorter100|7814_ ;
  assign \new_Sorter100|7915_  = \new_Sorter100|7815_  & \new_Sorter100|7816_ ;
  assign \new_Sorter100|7916_  = \new_Sorter100|7815_  | \new_Sorter100|7816_ ;
  assign \new_Sorter100|7917_  = \new_Sorter100|7817_  & \new_Sorter100|7818_ ;
  assign \new_Sorter100|7918_  = \new_Sorter100|7817_  | \new_Sorter100|7818_ ;
  assign \new_Sorter100|7919_  = \new_Sorter100|7819_  & \new_Sorter100|7820_ ;
  assign \new_Sorter100|7920_  = \new_Sorter100|7819_  | \new_Sorter100|7820_ ;
  assign \new_Sorter100|7921_  = \new_Sorter100|7821_  & \new_Sorter100|7822_ ;
  assign \new_Sorter100|7922_  = \new_Sorter100|7821_  | \new_Sorter100|7822_ ;
  assign \new_Sorter100|7923_  = \new_Sorter100|7823_  & \new_Sorter100|7824_ ;
  assign \new_Sorter100|7924_  = \new_Sorter100|7823_  | \new_Sorter100|7824_ ;
  assign \new_Sorter100|7925_  = \new_Sorter100|7825_  & \new_Sorter100|7826_ ;
  assign \new_Sorter100|7926_  = \new_Sorter100|7825_  | \new_Sorter100|7826_ ;
  assign \new_Sorter100|7927_  = \new_Sorter100|7827_  & \new_Sorter100|7828_ ;
  assign \new_Sorter100|7928_  = \new_Sorter100|7827_  | \new_Sorter100|7828_ ;
  assign \new_Sorter100|7929_  = \new_Sorter100|7829_  & \new_Sorter100|7830_ ;
  assign \new_Sorter100|7930_  = \new_Sorter100|7829_  | \new_Sorter100|7830_ ;
  assign \new_Sorter100|7931_  = \new_Sorter100|7831_  & \new_Sorter100|7832_ ;
  assign \new_Sorter100|7932_  = \new_Sorter100|7831_  | \new_Sorter100|7832_ ;
  assign \new_Sorter100|7933_  = \new_Sorter100|7833_  & \new_Sorter100|7834_ ;
  assign \new_Sorter100|7934_  = \new_Sorter100|7833_  | \new_Sorter100|7834_ ;
  assign \new_Sorter100|7935_  = \new_Sorter100|7835_  & \new_Sorter100|7836_ ;
  assign \new_Sorter100|7936_  = \new_Sorter100|7835_  | \new_Sorter100|7836_ ;
  assign \new_Sorter100|7937_  = \new_Sorter100|7837_  & \new_Sorter100|7838_ ;
  assign \new_Sorter100|7938_  = \new_Sorter100|7837_  | \new_Sorter100|7838_ ;
  assign \new_Sorter100|7939_  = \new_Sorter100|7839_  & \new_Sorter100|7840_ ;
  assign \new_Sorter100|7940_  = \new_Sorter100|7839_  | \new_Sorter100|7840_ ;
  assign \new_Sorter100|7941_  = \new_Sorter100|7841_  & \new_Sorter100|7842_ ;
  assign \new_Sorter100|7942_  = \new_Sorter100|7841_  | \new_Sorter100|7842_ ;
  assign \new_Sorter100|7943_  = \new_Sorter100|7843_  & \new_Sorter100|7844_ ;
  assign \new_Sorter100|7944_  = \new_Sorter100|7843_  | \new_Sorter100|7844_ ;
  assign \new_Sorter100|7945_  = \new_Sorter100|7845_  & \new_Sorter100|7846_ ;
  assign \new_Sorter100|7946_  = \new_Sorter100|7845_  | \new_Sorter100|7846_ ;
  assign \new_Sorter100|7947_  = \new_Sorter100|7847_  & \new_Sorter100|7848_ ;
  assign \new_Sorter100|7948_  = \new_Sorter100|7847_  | \new_Sorter100|7848_ ;
  assign \new_Sorter100|7949_  = \new_Sorter100|7849_  & \new_Sorter100|7850_ ;
  assign \new_Sorter100|7950_  = \new_Sorter100|7849_  | \new_Sorter100|7850_ ;
  assign \new_Sorter100|7951_  = \new_Sorter100|7851_  & \new_Sorter100|7852_ ;
  assign \new_Sorter100|7952_  = \new_Sorter100|7851_  | \new_Sorter100|7852_ ;
  assign \new_Sorter100|7953_  = \new_Sorter100|7853_  & \new_Sorter100|7854_ ;
  assign \new_Sorter100|7954_  = \new_Sorter100|7853_  | \new_Sorter100|7854_ ;
  assign \new_Sorter100|7955_  = \new_Sorter100|7855_  & \new_Sorter100|7856_ ;
  assign \new_Sorter100|7956_  = \new_Sorter100|7855_  | \new_Sorter100|7856_ ;
  assign \new_Sorter100|7957_  = \new_Sorter100|7857_  & \new_Sorter100|7858_ ;
  assign \new_Sorter100|7958_  = \new_Sorter100|7857_  | \new_Sorter100|7858_ ;
  assign \new_Sorter100|7959_  = \new_Sorter100|7859_  & \new_Sorter100|7860_ ;
  assign \new_Sorter100|7960_  = \new_Sorter100|7859_  | \new_Sorter100|7860_ ;
  assign \new_Sorter100|7961_  = \new_Sorter100|7861_  & \new_Sorter100|7862_ ;
  assign \new_Sorter100|7962_  = \new_Sorter100|7861_  | \new_Sorter100|7862_ ;
  assign \new_Sorter100|7963_  = \new_Sorter100|7863_  & \new_Sorter100|7864_ ;
  assign \new_Sorter100|7964_  = \new_Sorter100|7863_  | \new_Sorter100|7864_ ;
  assign \new_Sorter100|7965_  = \new_Sorter100|7865_  & \new_Sorter100|7866_ ;
  assign \new_Sorter100|7966_  = \new_Sorter100|7865_  | \new_Sorter100|7866_ ;
  assign \new_Sorter100|7967_  = \new_Sorter100|7867_  & \new_Sorter100|7868_ ;
  assign \new_Sorter100|7968_  = \new_Sorter100|7867_  | \new_Sorter100|7868_ ;
  assign \new_Sorter100|7969_  = \new_Sorter100|7869_  & \new_Sorter100|7870_ ;
  assign \new_Sorter100|7970_  = \new_Sorter100|7869_  | \new_Sorter100|7870_ ;
  assign \new_Sorter100|7971_  = \new_Sorter100|7871_  & \new_Sorter100|7872_ ;
  assign \new_Sorter100|7972_  = \new_Sorter100|7871_  | \new_Sorter100|7872_ ;
  assign \new_Sorter100|7973_  = \new_Sorter100|7873_  & \new_Sorter100|7874_ ;
  assign \new_Sorter100|7974_  = \new_Sorter100|7873_  | \new_Sorter100|7874_ ;
  assign \new_Sorter100|7975_  = \new_Sorter100|7875_  & \new_Sorter100|7876_ ;
  assign \new_Sorter100|7976_  = \new_Sorter100|7875_  | \new_Sorter100|7876_ ;
  assign \new_Sorter100|7977_  = \new_Sorter100|7877_  & \new_Sorter100|7878_ ;
  assign \new_Sorter100|7978_  = \new_Sorter100|7877_  | \new_Sorter100|7878_ ;
  assign \new_Sorter100|7979_  = \new_Sorter100|7879_  & \new_Sorter100|7880_ ;
  assign \new_Sorter100|7980_  = \new_Sorter100|7879_  | \new_Sorter100|7880_ ;
  assign \new_Sorter100|7981_  = \new_Sorter100|7881_  & \new_Sorter100|7882_ ;
  assign \new_Sorter100|7982_  = \new_Sorter100|7881_  | \new_Sorter100|7882_ ;
  assign \new_Sorter100|7983_  = \new_Sorter100|7883_  & \new_Sorter100|7884_ ;
  assign \new_Sorter100|7984_  = \new_Sorter100|7883_  | \new_Sorter100|7884_ ;
  assign \new_Sorter100|7985_  = \new_Sorter100|7885_  & \new_Sorter100|7886_ ;
  assign \new_Sorter100|7986_  = \new_Sorter100|7885_  | \new_Sorter100|7886_ ;
  assign \new_Sorter100|7987_  = \new_Sorter100|7887_  & \new_Sorter100|7888_ ;
  assign \new_Sorter100|7988_  = \new_Sorter100|7887_  | \new_Sorter100|7888_ ;
  assign \new_Sorter100|7989_  = \new_Sorter100|7889_  & \new_Sorter100|7890_ ;
  assign \new_Sorter100|7990_  = \new_Sorter100|7889_  | \new_Sorter100|7890_ ;
  assign \new_Sorter100|7991_  = \new_Sorter100|7891_  & \new_Sorter100|7892_ ;
  assign \new_Sorter100|7992_  = \new_Sorter100|7891_  | \new_Sorter100|7892_ ;
  assign \new_Sorter100|7993_  = \new_Sorter100|7893_  & \new_Sorter100|7894_ ;
  assign \new_Sorter100|7994_  = \new_Sorter100|7893_  | \new_Sorter100|7894_ ;
  assign \new_Sorter100|7995_  = \new_Sorter100|7895_  & \new_Sorter100|7896_ ;
  assign \new_Sorter100|7996_  = \new_Sorter100|7895_  | \new_Sorter100|7896_ ;
  assign \new_Sorter100|7997_  = \new_Sorter100|7897_  & \new_Sorter100|7898_ ;
  assign \new_Sorter100|7998_  = \new_Sorter100|7897_  | \new_Sorter100|7898_ ;
  assign \new_Sorter100|8000_  = \new_Sorter100|7900_  & \new_Sorter100|7901_ ;
  assign \new_Sorter100|8001_  = \new_Sorter100|7900_  | \new_Sorter100|7901_ ;
  assign \new_Sorter100|8002_  = \new_Sorter100|7902_  & \new_Sorter100|7903_ ;
  assign \new_Sorter100|8003_  = \new_Sorter100|7902_  | \new_Sorter100|7903_ ;
  assign \new_Sorter100|8004_  = \new_Sorter100|7904_  & \new_Sorter100|7905_ ;
  assign \new_Sorter100|8005_  = \new_Sorter100|7904_  | \new_Sorter100|7905_ ;
  assign \new_Sorter100|8006_  = \new_Sorter100|7906_  & \new_Sorter100|7907_ ;
  assign \new_Sorter100|8007_  = \new_Sorter100|7906_  | \new_Sorter100|7907_ ;
  assign \new_Sorter100|8008_  = \new_Sorter100|7908_  & \new_Sorter100|7909_ ;
  assign \new_Sorter100|8009_  = \new_Sorter100|7908_  | \new_Sorter100|7909_ ;
  assign \new_Sorter100|8010_  = \new_Sorter100|7910_  & \new_Sorter100|7911_ ;
  assign \new_Sorter100|8011_  = \new_Sorter100|7910_  | \new_Sorter100|7911_ ;
  assign \new_Sorter100|8012_  = \new_Sorter100|7912_  & \new_Sorter100|7913_ ;
  assign \new_Sorter100|8013_  = \new_Sorter100|7912_  | \new_Sorter100|7913_ ;
  assign \new_Sorter100|8014_  = \new_Sorter100|7914_  & \new_Sorter100|7915_ ;
  assign \new_Sorter100|8015_  = \new_Sorter100|7914_  | \new_Sorter100|7915_ ;
  assign \new_Sorter100|8016_  = \new_Sorter100|7916_  & \new_Sorter100|7917_ ;
  assign \new_Sorter100|8017_  = \new_Sorter100|7916_  | \new_Sorter100|7917_ ;
  assign \new_Sorter100|8018_  = \new_Sorter100|7918_  & \new_Sorter100|7919_ ;
  assign \new_Sorter100|8019_  = \new_Sorter100|7918_  | \new_Sorter100|7919_ ;
  assign \new_Sorter100|8020_  = \new_Sorter100|7920_  & \new_Sorter100|7921_ ;
  assign \new_Sorter100|8021_  = \new_Sorter100|7920_  | \new_Sorter100|7921_ ;
  assign \new_Sorter100|8022_  = \new_Sorter100|7922_  & \new_Sorter100|7923_ ;
  assign \new_Sorter100|8023_  = \new_Sorter100|7922_  | \new_Sorter100|7923_ ;
  assign \new_Sorter100|8024_  = \new_Sorter100|7924_  & \new_Sorter100|7925_ ;
  assign \new_Sorter100|8025_  = \new_Sorter100|7924_  | \new_Sorter100|7925_ ;
  assign \new_Sorter100|8026_  = \new_Sorter100|7926_  & \new_Sorter100|7927_ ;
  assign \new_Sorter100|8027_  = \new_Sorter100|7926_  | \new_Sorter100|7927_ ;
  assign \new_Sorter100|8028_  = \new_Sorter100|7928_  & \new_Sorter100|7929_ ;
  assign \new_Sorter100|8029_  = \new_Sorter100|7928_  | \new_Sorter100|7929_ ;
  assign \new_Sorter100|8030_  = \new_Sorter100|7930_  & \new_Sorter100|7931_ ;
  assign \new_Sorter100|8031_  = \new_Sorter100|7930_  | \new_Sorter100|7931_ ;
  assign \new_Sorter100|8032_  = \new_Sorter100|7932_  & \new_Sorter100|7933_ ;
  assign \new_Sorter100|8033_  = \new_Sorter100|7932_  | \new_Sorter100|7933_ ;
  assign \new_Sorter100|8034_  = \new_Sorter100|7934_  & \new_Sorter100|7935_ ;
  assign \new_Sorter100|8035_  = \new_Sorter100|7934_  | \new_Sorter100|7935_ ;
  assign \new_Sorter100|8036_  = \new_Sorter100|7936_  & \new_Sorter100|7937_ ;
  assign \new_Sorter100|8037_  = \new_Sorter100|7936_  | \new_Sorter100|7937_ ;
  assign \new_Sorter100|8038_  = \new_Sorter100|7938_  & \new_Sorter100|7939_ ;
  assign \new_Sorter100|8039_  = \new_Sorter100|7938_  | \new_Sorter100|7939_ ;
  assign \new_Sorter100|8040_  = \new_Sorter100|7940_  & \new_Sorter100|7941_ ;
  assign \new_Sorter100|8041_  = \new_Sorter100|7940_  | \new_Sorter100|7941_ ;
  assign \new_Sorter100|8042_  = \new_Sorter100|7942_  & \new_Sorter100|7943_ ;
  assign \new_Sorter100|8043_  = \new_Sorter100|7942_  | \new_Sorter100|7943_ ;
  assign \new_Sorter100|8044_  = \new_Sorter100|7944_  & \new_Sorter100|7945_ ;
  assign \new_Sorter100|8045_  = \new_Sorter100|7944_  | \new_Sorter100|7945_ ;
  assign \new_Sorter100|8046_  = \new_Sorter100|7946_  & \new_Sorter100|7947_ ;
  assign \new_Sorter100|8047_  = \new_Sorter100|7946_  | \new_Sorter100|7947_ ;
  assign \new_Sorter100|8048_  = \new_Sorter100|7948_  & \new_Sorter100|7949_ ;
  assign \new_Sorter100|8049_  = \new_Sorter100|7948_  | \new_Sorter100|7949_ ;
  assign \new_Sorter100|8050_  = \new_Sorter100|7950_  & \new_Sorter100|7951_ ;
  assign \new_Sorter100|8051_  = \new_Sorter100|7950_  | \new_Sorter100|7951_ ;
  assign \new_Sorter100|8052_  = \new_Sorter100|7952_  & \new_Sorter100|7953_ ;
  assign \new_Sorter100|8053_  = \new_Sorter100|7952_  | \new_Sorter100|7953_ ;
  assign \new_Sorter100|8054_  = \new_Sorter100|7954_  & \new_Sorter100|7955_ ;
  assign \new_Sorter100|8055_  = \new_Sorter100|7954_  | \new_Sorter100|7955_ ;
  assign \new_Sorter100|8056_  = \new_Sorter100|7956_  & \new_Sorter100|7957_ ;
  assign \new_Sorter100|8057_  = \new_Sorter100|7956_  | \new_Sorter100|7957_ ;
  assign \new_Sorter100|8058_  = \new_Sorter100|7958_  & \new_Sorter100|7959_ ;
  assign \new_Sorter100|8059_  = \new_Sorter100|7958_  | \new_Sorter100|7959_ ;
  assign \new_Sorter100|8060_  = \new_Sorter100|7960_  & \new_Sorter100|7961_ ;
  assign \new_Sorter100|8061_  = \new_Sorter100|7960_  | \new_Sorter100|7961_ ;
  assign \new_Sorter100|8062_  = \new_Sorter100|7962_  & \new_Sorter100|7963_ ;
  assign \new_Sorter100|8063_  = \new_Sorter100|7962_  | \new_Sorter100|7963_ ;
  assign \new_Sorter100|8064_  = \new_Sorter100|7964_  & \new_Sorter100|7965_ ;
  assign \new_Sorter100|8065_  = \new_Sorter100|7964_  | \new_Sorter100|7965_ ;
  assign \new_Sorter100|8066_  = \new_Sorter100|7966_  & \new_Sorter100|7967_ ;
  assign \new_Sorter100|8067_  = \new_Sorter100|7966_  | \new_Sorter100|7967_ ;
  assign \new_Sorter100|8068_  = \new_Sorter100|7968_  & \new_Sorter100|7969_ ;
  assign \new_Sorter100|8069_  = \new_Sorter100|7968_  | \new_Sorter100|7969_ ;
  assign \new_Sorter100|8070_  = \new_Sorter100|7970_  & \new_Sorter100|7971_ ;
  assign \new_Sorter100|8071_  = \new_Sorter100|7970_  | \new_Sorter100|7971_ ;
  assign \new_Sorter100|8072_  = \new_Sorter100|7972_  & \new_Sorter100|7973_ ;
  assign \new_Sorter100|8073_  = \new_Sorter100|7972_  | \new_Sorter100|7973_ ;
  assign \new_Sorter100|8074_  = \new_Sorter100|7974_  & \new_Sorter100|7975_ ;
  assign \new_Sorter100|8075_  = \new_Sorter100|7974_  | \new_Sorter100|7975_ ;
  assign \new_Sorter100|8076_  = \new_Sorter100|7976_  & \new_Sorter100|7977_ ;
  assign \new_Sorter100|8077_  = \new_Sorter100|7976_  | \new_Sorter100|7977_ ;
  assign \new_Sorter100|8078_  = \new_Sorter100|7978_  & \new_Sorter100|7979_ ;
  assign \new_Sorter100|8079_  = \new_Sorter100|7978_  | \new_Sorter100|7979_ ;
  assign \new_Sorter100|8080_  = \new_Sorter100|7980_  & \new_Sorter100|7981_ ;
  assign \new_Sorter100|8081_  = \new_Sorter100|7980_  | \new_Sorter100|7981_ ;
  assign \new_Sorter100|8082_  = \new_Sorter100|7982_  & \new_Sorter100|7983_ ;
  assign \new_Sorter100|8083_  = \new_Sorter100|7982_  | \new_Sorter100|7983_ ;
  assign \new_Sorter100|8084_  = \new_Sorter100|7984_  & \new_Sorter100|7985_ ;
  assign \new_Sorter100|8085_  = \new_Sorter100|7984_  | \new_Sorter100|7985_ ;
  assign \new_Sorter100|8086_  = \new_Sorter100|7986_  & \new_Sorter100|7987_ ;
  assign \new_Sorter100|8087_  = \new_Sorter100|7986_  | \new_Sorter100|7987_ ;
  assign \new_Sorter100|8088_  = \new_Sorter100|7988_  & \new_Sorter100|7989_ ;
  assign \new_Sorter100|8089_  = \new_Sorter100|7988_  | \new_Sorter100|7989_ ;
  assign \new_Sorter100|8090_  = \new_Sorter100|7990_  & \new_Sorter100|7991_ ;
  assign \new_Sorter100|8091_  = \new_Sorter100|7990_  | \new_Sorter100|7991_ ;
  assign \new_Sorter100|8092_  = \new_Sorter100|7992_  & \new_Sorter100|7993_ ;
  assign \new_Sorter100|8093_  = \new_Sorter100|7992_  | \new_Sorter100|7993_ ;
  assign \new_Sorter100|8094_  = \new_Sorter100|7994_  & \new_Sorter100|7995_ ;
  assign \new_Sorter100|8095_  = \new_Sorter100|7994_  | \new_Sorter100|7995_ ;
  assign \new_Sorter100|8096_  = \new_Sorter100|7996_  & \new_Sorter100|7997_ ;
  assign \new_Sorter100|8097_  = \new_Sorter100|7996_  | \new_Sorter100|7997_ ;
  assign \new_Sorter100|8098_  = \new_Sorter100|7998_  & \new_Sorter100|7999_ ;
  assign \new_Sorter100|8099_  = \new_Sorter100|7998_  | \new_Sorter100|7999_ ;
  assign \new_Sorter100|8100_  = \new_Sorter100|8000_ ;
  assign \new_Sorter100|8199_  = \new_Sorter100|8099_ ;
  assign \new_Sorter100|8101_  = \new_Sorter100|8001_  & \new_Sorter100|8002_ ;
  assign \new_Sorter100|8102_  = \new_Sorter100|8001_  | \new_Sorter100|8002_ ;
  assign \new_Sorter100|8103_  = \new_Sorter100|8003_  & \new_Sorter100|8004_ ;
  assign \new_Sorter100|8104_  = \new_Sorter100|8003_  | \new_Sorter100|8004_ ;
  assign \new_Sorter100|8105_  = \new_Sorter100|8005_  & \new_Sorter100|8006_ ;
  assign \new_Sorter100|8106_  = \new_Sorter100|8005_  | \new_Sorter100|8006_ ;
  assign \new_Sorter100|8107_  = \new_Sorter100|8007_  & \new_Sorter100|8008_ ;
  assign \new_Sorter100|8108_  = \new_Sorter100|8007_  | \new_Sorter100|8008_ ;
  assign \new_Sorter100|8109_  = \new_Sorter100|8009_  & \new_Sorter100|8010_ ;
  assign \new_Sorter100|8110_  = \new_Sorter100|8009_  | \new_Sorter100|8010_ ;
  assign \new_Sorter100|8111_  = \new_Sorter100|8011_  & \new_Sorter100|8012_ ;
  assign \new_Sorter100|8112_  = \new_Sorter100|8011_  | \new_Sorter100|8012_ ;
  assign \new_Sorter100|8113_  = \new_Sorter100|8013_  & \new_Sorter100|8014_ ;
  assign \new_Sorter100|8114_  = \new_Sorter100|8013_  | \new_Sorter100|8014_ ;
  assign \new_Sorter100|8115_  = \new_Sorter100|8015_  & \new_Sorter100|8016_ ;
  assign \new_Sorter100|8116_  = \new_Sorter100|8015_  | \new_Sorter100|8016_ ;
  assign \new_Sorter100|8117_  = \new_Sorter100|8017_  & \new_Sorter100|8018_ ;
  assign \new_Sorter100|8118_  = \new_Sorter100|8017_  | \new_Sorter100|8018_ ;
  assign \new_Sorter100|8119_  = \new_Sorter100|8019_  & \new_Sorter100|8020_ ;
  assign \new_Sorter100|8120_  = \new_Sorter100|8019_  | \new_Sorter100|8020_ ;
  assign \new_Sorter100|8121_  = \new_Sorter100|8021_  & \new_Sorter100|8022_ ;
  assign \new_Sorter100|8122_  = \new_Sorter100|8021_  | \new_Sorter100|8022_ ;
  assign \new_Sorter100|8123_  = \new_Sorter100|8023_  & \new_Sorter100|8024_ ;
  assign \new_Sorter100|8124_  = \new_Sorter100|8023_  | \new_Sorter100|8024_ ;
  assign \new_Sorter100|8125_  = \new_Sorter100|8025_  & \new_Sorter100|8026_ ;
  assign \new_Sorter100|8126_  = \new_Sorter100|8025_  | \new_Sorter100|8026_ ;
  assign \new_Sorter100|8127_  = \new_Sorter100|8027_  & \new_Sorter100|8028_ ;
  assign \new_Sorter100|8128_  = \new_Sorter100|8027_  | \new_Sorter100|8028_ ;
  assign \new_Sorter100|8129_  = \new_Sorter100|8029_  & \new_Sorter100|8030_ ;
  assign \new_Sorter100|8130_  = \new_Sorter100|8029_  | \new_Sorter100|8030_ ;
  assign \new_Sorter100|8131_  = \new_Sorter100|8031_  & \new_Sorter100|8032_ ;
  assign \new_Sorter100|8132_  = \new_Sorter100|8031_  | \new_Sorter100|8032_ ;
  assign \new_Sorter100|8133_  = \new_Sorter100|8033_  & \new_Sorter100|8034_ ;
  assign \new_Sorter100|8134_  = \new_Sorter100|8033_  | \new_Sorter100|8034_ ;
  assign \new_Sorter100|8135_  = \new_Sorter100|8035_  & \new_Sorter100|8036_ ;
  assign \new_Sorter100|8136_  = \new_Sorter100|8035_  | \new_Sorter100|8036_ ;
  assign \new_Sorter100|8137_  = \new_Sorter100|8037_  & \new_Sorter100|8038_ ;
  assign \new_Sorter100|8138_  = \new_Sorter100|8037_  | \new_Sorter100|8038_ ;
  assign \new_Sorter100|8139_  = \new_Sorter100|8039_  & \new_Sorter100|8040_ ;
  assign \new_Sorter100|8140_  = \new_Sorter100|8039_  | \new_Sorter100|8040_ ;
  assign \new_Sorter100|8141_  = \new_Sorter100|8041_  & \new_Sorter100|8042_ ;
  assign \new_Sorter100|8142_  = \new_Sorter100|8041_  | \new_Sorter100|8042_ ;
  assign \new_Sorter100|8143_  = \new_Sorter100|8043_  & \new_Sorter100|8044_ ;
  assign \new_Sorter100|8144_  = \new_Sorter100|8043_  | \new_Sorter100|8044_ ;
  assign \new_Sorter100|8145_  = \new_Sorter100|8045_  & \new_Sorter100|8046_ ;
  assign \new_Sorter100|8146_  = \new_Sorter100|8045_  | \new_Sorter100|8046_ ;
  assign \new_Sorter100|8147_  = \new_Sorter100|8047_  & \new_Sorter100|8048_ ;
  assign \new_Sorter100|8148_  = \new_Sorter100|8047_  | \new_Sorter100|8048_ ;
  assign \new_Sorter100|8149_  = \new_Sorter100|8049_  & \new_Sorter100|8050_ ;
  assign \new_Sorter100|8150_  = \new_Sorter100|8049_  | \new_Sorter100|8050_ ;
  assign \new_Sorter100|8151_  = \new_Sorter100|8051_  & \new_Sorter100|8052_ ;
  assign \new_Sorter100|8152_  = \new_Sorter100|8051_  | \new_Sorter100|8052_ ;
  assign \new_Sorter100|8153_  = \new_Sorter100|8053_  & \new_Sorter100|8054_ ;
  assign \new_Sorter100|8154_  = \new_Sorter100|8053_  | \new_Sorter100|8054_ ;
  assign \new_Sorter100|8155_  = \new_Sorter100|8055_  & \new_Sorter100|8056_ ;
  assign \new_Sorter100|8156_  = \new_Sorter100|8055_  | \new_Sorter100|8056_ ;
  assign \new_Sorter100|8157_  = \new_Sorter100|8057_  & \new_Sorter100|8058_ ;
  assign \new_Sorter100|8158_  = \new_Sorter100|8057_  | \new_Sorter100|8058_ ;
  assign \new_Sorter100|8159_  = \new_Sorter100|8059_  & \new_Sorter100|8060_ ;
  assign \new_Sorter100|8160_  = \new_Sorter100|8059_  | \new_Sorter100|8060_ ;
  assign \new_Sorter100|8161_  = \new_Sorter100|8061_  & \new_Sorter100|8062_ ;
  assign \new_Sorter100|8162_  = \new_Sorter100|8061_  | \new_Sorter100|8062_ ;
  assign \new_Sorter100|8163_  = \new_Sorter100|8063_  & \new_Sorter100|8064_ ;
  assign \new_Sorter100|8164_  = \new_Sorter100|8063_  | \new_Sorter100|8064_ ;
  assign \new_Sorter100|8165_  = \new_Sorter100|8065_  & \new_Sorter100|8066_ ;
  assign \new_Sorter100|8166_  = \new_Sorter100|8065_  | \new_Sorter100|8066_ ;
  assign \new_Sorter100|8167_  = \new_Sorter100|8067_  & \new_Sorter100|8068_ ;
  assign \new_Sorter100|8168_  = \new_Sorter100|8067_  | \new_Sorter100|8068_ ;
  assign \new_Sorter100|8169_  = \new_Sorter100|8069_  & \new_Sorter100|8070_ ;
  assign \new_Sorter100|8170_  = \new_Sorter100|8069_  | \new_Sorter100|8070_ ;
  assign \new_Sorter100|8171_  = \new_Sorter100|8071_  & \new_Sorter100|8072_ ;
  assign \new_Sorter100|8172_  = \new_Sorter100|8071_  | \new_Sorter100|8072_ ;
  assign \new_Sorter100|8173_  = \new_Sorter100|8073_  & \new_Sorter100|8074_ ;
  assign \new_Sorter100|8174_  = \new_Sorter100|8073_  | \new_Sorter100|8074_ ;
  assign \new_Sorter100|8175_  = \new_Sorter100|8075_  & \new_Sorter100|8076_ ;
  assign \new_Sorter100|8176_  = \new_Sorter100|8075_  | \new_Sorter100|8076_ ;
  assign \new_Sorter100|8177_  = \new_Sorter100|8077_  & \new_Sorter100|8078_ ;
  assign \new_Sorter100|8178_  = \new_Sorter100|8077_  | \new_Sorter100|8078_ ;
  assign \new_Sorter100|8179_  = \new_Sorter100|8079_  & \new_Sorter100|8080_ ;
  assign \new_Sorter100|8180_  = \new_Sorter100|8079_  | \new_Sorter100|8080_ ;
  assign \new_Sorter100|8181_  = \new_Sorter100|8081_  & \new_Sorter100|8082_ ;
  assign \new_Sorter100|8182_  = \new_Sorter100|8081_  | \new_Sorter100|8082_ ;
  assign \new_Sorter100|8183_  = \new_Sorter100|8083_  & \new_Sorter100|8084_ ;
  assign \new_Sorter100|8184_  = \new_Sorter100|8083_  | \new_Sorter100|8084_ ;
  assign \new_Sorter100|8185_  = \new_Sorter100|8085_  & \new_Sorter100|8086_ ;
  assign \new_Sorter100|8186_  = \new_Sorter100|8085_  | \new_Sorter100|8086_ ;
  assign \new_Sorter100|8187_  = \new_Sorter100|8087_  & \new_Sorter100|8088_ ;
  assign \new_Sorter100|8188_  = \new_Sorter100|8087_  | \new_Sorter100|8088_ ;
  assign \new_Sorter100|8189_  = \new_Sorter100|8089_  & \new_Sorter100|8090_ ;
  assign \new_Sorter100|8190_  = \new_Sorter100|8089_  | \new_Sorter100|8090_ ;
  assign \new_Sorter100|8191_  = \new_Sorter100|8091_  & \new_Sorter100|8092_ ;
  assign \new_Sorter100|8192_  = \new_Sorter100|8091_  | \new_Sorter100|8092_ ;
  assign \new_Sorter100|8193_  = \new_Sorter100|8093_  & \new_Sorter100|8094_ ;
  assign \new_Sorter100|8194_  = \new_Sorter100|8093_  | \new_Sorter100|8094_ ;
  assign \new_Sorter100|8195_  = \new_Sorter100|8095_  & \new_Sorter100|8096_ ;
  assign \new_Sorter100|8196_  = \new_Sorter100|8095_  | \new_Sorter100|8096_ ;
  assign \new_Sorter100|8197_  = \new_Sorter100|8097_  & \new_Sorter100|8098_ ;
  assign \new_Sorter100|8198_  = \new_Sorter100|8097_  | \new_Sorter100|8098_ ;
  assign \new_Sorter100|8200_  = \new_Sorter100|8100_  & \new_Sorter100|8101_ ;
  assign \new_Sorter100|8201_  = \new_Sorter100|8100_  | \new_Sorter100|8101_ ;
  assign \new_Sorter100|8202_  = \new_Sorter100|8102_  & \new_Sorter100|8103_ ;
  assign \new_Sorter100|8203_  = \new_Sorter100|8102_  | \new_Sorter100|8103_ ;
  assign \new_Sorter100|8204_  = \new_Sorter100|8104_  & \new_Sorter100|8105_ ;
  assign \new_Sorter100|8205_  = \new_Sorter100|8104_  | \new_Sorter100|8105_ ;
  assign \new_Sorter100|8206_  = \new_Sorter100|8106_  & \new_Sorter100|8107_ ;
  assign \new_Sorter100|8207_  = \new_Sorter100|8106_  | \new_Sorter100|8107_ ;
  assign \new_Sorter100|8208_  = \new_Sorter100|8108_  & \new_Sorter100|8109_ ;
  assign \new_Sorter100|8209_  = \new_Sorter100|8108_  | \new_Sorter100|8109_ ;
  assign \new_Sorter100|8210_  = \new_Sorter100|8110_  & \new_Sorter100|8111_ ;
  assign \new_Sorter100|8211_  = \new_Sorter100|8110_  | \new_Sorter100|8111_ ;
  assign \new_Sorter100|8212_  = \new_Sorter100|8112_  & \new_Sorter100|8113_ ;
  assign \new_Sorter100|8213_  = \new_Sorter100|8112_  | \new_Sorter100|8113_ ;
  assign \new_Sorter100|8214_  = \new_Sorter100|8114_  & \new_Sorter100|8115_ ;
  assign \new_Sorter100|8215_  = \new_Sorter100|8114_  | \new_Sorter100|8115_ ;
  assign \new_Sorter100|8216_  = \new_Sorter100|8116_  & \new_Sorter100|8117_ ;
  assign \new_Sorter100|8217_  = \new_Sorter100|8116_  | \new_Sorter100|8117_ ;
  assign \new_Sorter100|8218_  = \new_Sorter100|8118_  & \new_Sorter100|8119_ ;
  assign \new_Sorter100|8219_  = \new_Sorter100|8118_  | \new_Sorter100|8119_ ;
  assign \new_Sorter100|8220_  = \new_Sorter100|8120_  & \new_Sorter100|8121_ ;
  assign \new_Sorter100|8221_  = \new_Sorter100|8120_  | \new_Sorter100|8121_ ;
  assign \new_Sorter100|8222_  = \new_Sorter100|8122_  & \new_Sorter100|8123_ ;
  assign \new_Sorter100|8223_  = \new_Sorter100|8122_  | \new_Sorter100|8123_ ;
  assign \new_Sorter100|8224_  = \new_Sorter100|8124_  & \new_Sorter100|8125_ ;
  assign \new_Sorter100|8225_  = \new_Sorter100|8124_  | \new_Sorter100|8125_ ;
  assign \new_Sorter100|8226_  = \new_Sorter100|8126_  & \new_Sorter100|8127_ ;
  assign \new_Sorter100|8227_  = \new_Sorter100|8126_  | \new_Sorter100|8127_ ;
  assign \new_Sorter100|8228_  = \new_Sorter100|8128_  & \new_Sorter100|8129_ ;
  assign \new_Sorter100|8229_  = \new_Sorter100|8128_  | \new_Sorter100|8129_ ;
  assign \new_Sorter100|8230_  = \new_Sorter100|8130_  & \new_Sorter100|8131_ ;
  assign \new_Sorter100|8231_  = \new_Sorter100|8130_  | \new_Sorter100|8131_ ;
  assign \new_Sorter100|8232_  = \new_Sorter100|8132_  & \new_Sorter100|8133_ ;
  assign \new_Sorter100|8233_  = \new_Sorter100|8132_  | \new_Sorter100|8133_ ;
  assign \new_Sorter100|8234_  = \new_Sorter100|8134_  & \new_Sorter100|8135_ ;
  assign \new_Sorter100|8235_  = \new_Sorter100|8134_  | \new_Sorter100|8135_ ;
  assign \new_Sorter100|8236_  = \new_Sorter100|8136_  & \new_Sorter100|8137_ ;
  assign \new_Sorter100|8237_  = \new_Sorter100|8136_  | \new_Sorter100|8137_ ;
  assign \new_Sorter100|8238_  = \new_Sorter100|8138_  & \new_Sorter100|8139_ ;
  assign \new_Sorter100|8239_  = \new_Sorter100|8138_  | \new_Sorter100|8139_ ;
  assign \new_Sorter100|8240_  = \new_Sorter100|8140_  & \new_Sorter100|8141_ ;
  assign \new_Sorter100|8241_  = \new_Sorter100|8140_  | \new_Sorter100|8141_ ;
  assign \new_Sorter100|8242_  = \new_Sorter100|8142_  & \new_Sorter100|8143_ ;
  assign \new_Sorter100|8243_  = \new_Sorter100|8142_  | \new_Sorter100|8143_ ;
  assign \new_Sorter100|8244_  = \new_Sorter100|8144_  & \new_Sorter100|8145_ ;
  assign \new_Sorter100|8245_  = \new_Sorter100|8144_  | \new_Sorter100|8145_ ;
  assign \new_Sorter100|8246_  = \new_Sorter100|8146_  & \new_Sorter100|8147_ ;
  assign \new_Sorter100|8247_  = \new_Sorter100|8146_  | \new_Sorter100|8147_ ;
  assign \new_Sorter100|8248_  = \new_Sorter100|8148_  & \new_Sorter100|8149_ ;
  assign \new_Sorter100|8249_  = \new_Sorter100|8148_  | \new_Sorter100|8149_ ;
  assign \new_Sorter100|8250_  = \new_Sorter100|8150_  & \new_Sorter100|8151_ ;
  assign \new_Sorter100|8251_  = \new_Sorter100|8150_  | \new_Sorter100|8151_ ;
  assign \new_Sorter100|8252_  = \new_Sorter100|8152_  & \new_Sorter100|8153_ ;
  assign \new_Sorter100|8253_  = \new_Sorter100|8152_  | \new_Sorter100|8153_ ;
  assign \new_Sorter100|8254_  = \new_Sorter100|8154_  & \new_Sorter100|8155_ ;
  assign \new_Sorter100|8255_  = \new_Sorter100|8154_  | \new_Sorter100|8155_ ;
  assign \new_Sorter100|8256_  = \new_Sorter100|8156_  & \new_Sorter100|8157_ ;
  assign \new_Sorter100|8257_  = \new_Sorter100|8156_  | \new_Sorter100|8157_ ;
  assign \new_Sorter100|8258_  = \new_Sorter100|8158_  & \new_Sorter100|8159_ ;
  assign \new_Sorter100|8259_  = \new_Sorter100|8158_  | \new_Sorter100|8159_ ;
  assign \new_Sorter100|8260_  = \new_Sorter100|8160_  & \new_Sorter100|8161_ ;
  assign \new_Sorter100|8261_  = \new_Sorter100|8160_  | \new_Sorter100|8161_ ;
  assign \new_Sorter100|8262_  = \new_Sorter100|8162_  & \new_Sorter100|8163_ ;
  assign \new_Sorter100|8263_  = \new_Sorter100|8162_  | \new_Sorter100|8163_ ;
  assign \new_Sorter100|8264_  = \new_Sorter100|8164_  & \new_Sorter100|8165_ ;
  assign \new_Sorter100|8265_  = \new_Sorter100|8164_  | \new_Sorter100|8165_ ;
  assign \new_Sorter100|8266_  = \new_Sorter100|8166_  & \new_Sorter100|8167_ ;
  assign \new_Sorter100|8267_  = \new_Sorter100|8166_  | \new_Sorter100|8167_ ;
  assign \new_Sorter100|8268_  = \new_Sorter100|8168_  & \new_Sorter100|8169_ ;
  assign \new_Sorter100|8269_  = \new_Sorter100|8168_  | \new_Sorter100|8169_ ;
  assign \new_Sorter100|8270_  = \new_Sorter100|8170_  & \new_Sorter100|8171_ ;
  assign \new_Sorter100|8271_  = \new_Sorter100|8170_  | \new_Sorter100|8171_ ;
  assign \new_Sorter100|8272_  = \new_Sorter100|8172_  & \new_Sorter100|8173_ ;
  assign \new_Sorter100|8273_  = \new_Sorter100|8172_  | \new_Sorter100|8173_ ;
  assign \new_Sorter100|8274_  = \new_Sorter100|8174_  & \new_Sorter100|8175_ ;
  assign \new_Sorter100|8275_  = \new_Sorter100|8174_  | \new_Sorter100|8175_ ;
  assign \new_Sorter100|8276_  = \new_Sorter100|8176_  & \new_Sorter100|8177_ ;
  assign \new_Sorter100|8277_  = \new_Sorter100|8176_  | \new_Sorter100|8177_ ;
  assign \new_Sorter100|8278_  = \new_Sorter100|8178_  & \new_Sorter100|8179_ ;
  assign \new_Sorter100|8279_  = \new_Sorter100|8178_  | \new_Sorter100|8179_ ;
  assign \new_Sorter100|8280_  = \new_Sorter100|8180_  & \new_Sorter100|8181_ ;
  assign \new_Sorter100|8281_  = \new_Sorter100|8180_  | \new_Sorter100|8181_ ;
  assign \new_Sorter100|8282_  = \new_Sorter100|8182_  & \new_Sorter100|8183_ ;
  assign \new_Sorter100|8283_  = \new_Sorter100|8182_  | \new_Sorter100|8183_ ;
  assign \new_Sorter100|8284_  = \new_Sorter100|8184_  & \new_Sorter100|8185_ ;
  assign \new_Sorter100|8285_  = \new_Sorter100|8184_  | \new_Sorter100|8185_ ;
  assign \new_Sorter100|8286_  = \new_Sorter100|8186_  & \new_Sorter100|8187_ ;
  assign \new_Sorter100|8287_  = \new_Sorter100|8186_  | \new_Sorter100|8187_ ;
  assign \new_Sorter100|8288_  = \new_Sorter100|8188_  & \new_Sorter100|8189_ ;
  assign \new_Sorter100|8289_  = \new_Sorter100|8188_  | \new_Sorter100|8189_ ;
  assign \new_Sorter100|8290_  = \new_Sorter100|8190_  & \new_Sorter100|8191_ ;
  assign \new_Sorter100|8291_  = \new_Sorter100|8190_  | \new_Sorter100|8191_ ;
  assign \new_Sorter100|8292_  = \new_Sorter100|8192_  & \new_Sorter100|8193_ ;
  assign \new_Sorter100|8293_  = \new_Sorter100|8192_  | \new_Sorter100|8193_ ;
  assign \new_Sorter100|8294_  = \new_Sorter100|8194_  & \new_Sorter100|8195_ ;
  assign \new_Sorter100|8295_  = \new_Sorter100|8194_  | \new_Sorter100|8195_ ;
  assign \new_Sorter100|8296_  = \new_Sorter100|8196_  & \new_Sorter100|8197_ ;
  assign \new_Sorter100|8297_  = \new_Sorter100|8196_  | \new_Sorter100|8197_ ;
  assign \new_Sorter100|8298_  = \new_Sorter100|8198_  & \new_Sorter100|8199_ ;
  assign \new_Sorter100|8299_  = \new_Sorter100|8198_  | \new_Sorter100|8199_ ;
  assign \new_Sorter100|8300_  = \new_Sorter100|8200_ ;
  assign \new_Sorter100|8399_  = \new_Sorter100|8299_ ;
  assign \new_Sorter100|8301_  = \new_Sorter100|8201_  & \new_Sorter100|8202_ ;
  assign \new_Sorter100|8302_  = \new_Sorter100|8201_  | \new_Sorter100|8202_ ;
  assign \new_Sorter100|8303_  = \new_Sorter100|8203_  & \new_Sorter100|8204_ ;
  assign \new_Sorter100|8304_  = \new_Sorter100|8203_  | \new_Sorter100|8204_ ;
  assign \new_Sorter100|8305_  = \new_Sorter100|8205_  & \new_Sorter100|8206_ ;
  assign \new_Sorter100|8306_  = \new_Sorter100|8205_  | \new_Sorter100|8206_ ;
  assign \new_Sorter100|8307_  = \new_Sorter100|8207_  & \new_Sorter100|8208_ ;
  assign \new_Sorter100|8308_  = \new_Sorter100|8207_  | \new_Sorter100|8208_ ;
  assign \new_Sorter100|8309_  = \new_Sorter100|8209_  & \new_Sorter100|8210_ ;
  assign \new_Sorter100|8310_  = \new_Sorter100|8209_  | \new_Sorter100|8210_ ;
  assign \new_Sorter100|8311_  = \new_Sorter100|8211_  & \new_Sorter100|8212_ ;
  assign \new_Sorter100|8312_  = \new_Sorter100|8211_  | \new_Sorter100|8212_ ;
  assign \new_Sorter100|8313_  = \new_Sorter100|8213_  & \new_Sorter100|8214_ ;
  assign \new_Sorter100|8314_  = \new_Sorter100|8213_  | \new_Sorter100|8214_ ;
  assign \new_Sorter100|8315_  = \new_Sorter100|8215_  & \new_Sorter100|8216_ ;
  assign \new_Sorter100|8316_  = \new_Sorter100|8215_  | \new_Sorter100|8216_ ;
  assign \new_Sorter100|8317_  = \new_Sorter100|8217_  & \new_Sorter100|8218_ ;
  assign \new_Sorter100|8318_  = \new_Sorter100|8217_  | \new_Sorter100|8218_ ;
  assign \new_Sorter100|8319_  = \new_Sorter100|8219_  & \new_Sorter100|8220_ ;
  assign \new_Sorter100|8320_  = \new_Sorter100|8219_  | \new_Sorter100|8220_ ;
  assign \new_Sorter100|8321_  = \new_Sorter100|8221_  & \new_Sorter100|8222_ ;
  assign \new_Sorter100|8322_  = \new_Sorter100|8221_  | \new_Sorter100|8222_ ;
  assign \new_Sorter100|8323_  = \new_Sorter100|8223_  & \new_Sorter100|8224_ ;
  assign \new_Sorter100|8324_  = \new_Sorter100|8223_  | \new_Sorter100|8224_ ;
  assign \new_Sorter100|8325_  = \new_Sorter100|8225_  & \new_Sorter100|8226_ ;
  assign \new_Sorter100|8326_  = \new_Sorter100|8225_  | \new_Sorter100|8226_ ;
  assign \new_Sorter100|8327_  = \new_Sorter100|8227_  & \new_Sorter100|8228_ ;
  assign \new_Sorter100|8328_  = \new_Sorter100|8227_  | \new_Sorter100|8228_ ;
  assign \new_Sorter100|8329_  = \new_Sorter100|8229_  & \new_Sorter100|8230_ ;
  assign \new_Sorter100|8330_  = \new_Sorter100|8229_  | \new_Sorter100|8230_ ;
  assign \new_Sorter100|8331_  = \new_Sorter100|8231_  & \new_Sorter100|8232_ ;
  assign \new_Sorter100|8332_  = \new_Sorter100|8231_  | \new_Sorter100|8232_ ;
  assign \new_Sorter100|8333_  = \new_Sorter100|8233_  & \new_Sorter100|8234_ ;
  assign \new_Sorter100|8334_  = \new_Sorter100|8233_  | \new_Sorter100|8234_ ;
  assign \new_Sorter100|8335_  = \new_Sorter100|8235_  & \new_Sorter100|8236_ ;
  assign \new_Sorter100|8336_  = \new_Sorter100|8235_  | \new_Sorter100|8236_ ;
  assign \new_Sorter100|8337_  = \new_Sorter100|8237_  & \new_Sorter100|8238_ ;
  assign \new_Sorter100|8338_  = \new_Sorter100|8237_  | \new_Sorter100|8238_ ;
  assign \new_Sorter100|8339_  = \new_Sorter100|8239_  & \new_Sorter100|8240_ ;
  assign \new_Sorter100|8340_  = \new_Sorter100|8239_  | \new_Sorter100|8240_ ;
  assign \new_Sorter100|8341_  = \new_Sorter100|8241_  & \new_Sorter100|8242_ ;
  assign \new_Sorter100|8342_  = \new_Sorter100|8241_  | \new_Sorter100|8242_ ;
  assign \new_Sorter100|8343_  = \new_Sorter100|8243_  & \new_Sorter100|8244_ ;
  assign \new_Sorter100|8344_  = \new_Sorter100|8243_  | \new_Sorter100|8244_ ;
  assign \new_Sorter100|8345_  = \new_Sorter100|8245_  & \new_Sorter100|8246_ ;
  assign \new_Sorter100|8346_  = \new_Sorter100|8245_  | \new_Sorter100|8246_ ;
  assign \new_Sorter100|8347_  = \new_Sorter100|8247_  & \new_Sorter100|8248_ ;
  assign \new_Sorter100|8348_  = \new_Sorter100|8247_  | \new_Sorter100|8248_ ;
  assign \new_Sorter100|8349_  = \new_Sorter100|8249_  & \new_Sorter100|8250_ ;
  assign \new_Sorter100|8350_  = \new_Sorter100|8249_  | \new_Sorter100|8250_ ;
  assign \new_Sorter100|8351_  = \new_Sorter100|8251_  & \new_Sorter100|8252_ ;
  assign \new_Sorter100|8352_  = \new_Sorter100|8251_  | \new_Sorter100|8252_ ;
  assign \new_Sorter100|8353_  = \new_Sorter100|8253_  & \new_Sorter100|8254_ ;
  assign \new_Sorter100|8354_  = \new_Sorter100|8253_  | \new_Sorter100|8254_ ;
  assign \new_Sorter100|8355_  = \new_Sorter100|8255_  & \new_Sorter100|8256_ ;
  assign \new_Sorter100|8356_  = \new_Sorter100|8255_  | \new_Sorter100|8256_ ;
  assign \new_Sorter100|8357_  = \new_Sorter100|8257_  & \new_Sorter100|8258_ ;
  assign \new_Sorter100|8358_  = \new_Sorter100|8257_  | \new_Sorter100|8258_ ;
  assign \new_Sorter100|8359_  = \new_Sorter100|8259_  & \new_Sorter100|8260_ ;
  assign \new_Sorter100|8360_  = \new_Sorter100|8259_  | \new_Sorter100|8260_ ;
  assign \new_Sorter100|8361_  = \new_Sorter100|8261_  & \new_Sorter100|8262_ ;
  assign \new_Sorter100|8362_  = \new_Sorter100|8261_  | \new_Sorter100|8262_ ;
  assign \new_Sorter100|8363_  = \new_Sorter100|8263_  & \new_Sorter100|8264_ ;
  assign \new_Sorter100|8364_  = \new_Sorter100|8263_  | \new_Sorter100|8264_ ;
  assign \new_Sorter100|8365_  = \new_Sorter100|8265_  & \new_Sorter100|8266_ ;
  assign \new_Sorter100|8366_  = \new_Sorter100|8265_  | \new_Sorter100|8266_ ;
  assign \new_Sorter100|8367_  = \new_Sorter100|8267_  & \new_Sorter100|8268_ ;
  assign \new_Sorter100|8368_  = \new_Sorter100|8267_  | \new_Sorter100|8268_ ;
  assign \new_Sorter100|8369_  = \new_Sorter100|8269_  & \new_Sorter100|8270_ ;
  assign \new_Sorter100|8370_  = \new_Sorter100|8269_  | \new_Sorter100|8270_ ;
  assign \new_Sorter100|8371_  = \new_Sorter100|8271_  & \new_Sorter100|8272_ ;
  assign \new_Sorter100|8372_  = \new_Sorter100|8271_  | \new_Sorter100|8272_ ;
  assign \new_Sorter100|8373_  = \new_Sorter100|8273_  & \new_Sorter100|8274_ ;
  assign \new_Sorter100|8374_  = \new_Sorter100|8273_  | \new_Sorter100|8274_ ;
  assign \new_Sorter100|8375_  = \new_Sorter100|8275_  & \new_Sorter100|8276_ ;
  assign \new_Sorter100|8376_  = \new_Sorter100|8275_  | \new_Sorter100|8276_ ;
  assign \new_Sorter100|8377_  = \new_Sorter100|8277_  & \new_Sorter100|8278_ ;
  assign \new_Sorter100|8378_  = \new_Sorter100|8277_  | \new_Sorter100|8278_ ;
  assign \new_Sorter100|8379_  = \new_Sorter100|8279_  & \new_Sorter100|8280_ ;
  assign \new_Sorter100|8380_  = \new_Sorter100|8279_  | \new_Sorter100|8280_ ;
  assign \new_Sorter100|8381_  = \new_Sorter100|8281_  & \new_Sorter100|8282_ ;
  assign \new_Sorter100|8382_  = \new_Sorter100|8281_  | \new_Sorter100|8282_ ;
  assign \new_Sorter100|8383_  = \new_Sorter100|8283_  & \new_Sorter100|8284_ ;
  assign \new_Sorter100|8384_  = \new_Sorter100|8283_  | \new_Sorter100|8284_ ;
  assign \new_Sorter100|8385_  = \new_Sorter100|8285_  & \new_Sorter100|8286_ ;
  assign \new_Sorter100|8386_  = \new_Sorter100|8285_  | \new_Sorter100|8286_ ;
  assign \new_Sorter100|8387_  = \new_Sorter100|8287_  & \new_Sorter100|8288_ ;
  assign \new_Sorter100|8388_  = \new_Sorter100|8287_  | \new_Sorter100|8288_ ;
  assign \new_Sorter100|8389_  = \new_Sorter100|8289_  & \new_Sorter100|8290_ ;
  assign \new_Sorter100|8390_  = \new_Sorter100|8289_  | \new_Sorter100|8290_ ;
  assign \new_Sorter100|8391_  = \new_Sorter100|8291_  & \new_Sorter100|8292_ ;
  assign \new_Sorter100|8392_  = \new_Sorter100|8291_  | \new_Sorter100|8292_ ;
  assign \new_Sorter100|8393_  = \new_Sorter100|8293_  & \new_Sorter100|8294_ ;
  assign \new_Sorter100|8394_  = \new_Sorter100|8293_  | \new_Sorter100|8294_ ;
  assign \new_Sorter100|8395_  = \new_Sorter100|8295_  & \new_Sorter100|8296_ ;
  assign \new_Sorter100|8396_  = \new_Sorter100|8295_  | \new_Sorter100|8296_ ;
  assign \new_Sorter100|8397_  = \new_Sorter100|8297_  & \new_Sorter100|8298_ ;
  assign \new_Sorter100|8398_  = \new_Sorter100|8297_  | \new_Sorter100|8298_ ;
  assign \new_Sorter100|8400_  = \new_Sorter100|8300_  & \new_Sorter100|8301_ ;
  assign \new_Sorter100|8401_  = \new_Sorter100|8300_  | \new_Sorter100|8301_ ;
  assign \new_Sorter100|8402_  = \new_Sorter100|8302_  & \new_Sorter100|8303_ ;
  assign \new_Sorter100|8403_  = \new_Sorter100|8302_  | \new_Sorter100|8303_ ;
  assign \new_Sorter100|8404_  = \new_Sorter100|8304_  & \new_Sorter100|8305_ ;
  assign \new_Sorter100|8405_  = \new_Sorter100|8304_  | \new_Sorter100|8305_ ;
  assign \new_Sorter100|8406_  = \new_Sorter100|8306_  & \new_Sorter100|8307_ ;
  assign \new_Sorter100|8407_  = \new_Sorter100|8306_  | \new_Sorter100|8307_ ;
  assign \new_Sorter100|8408_  = \new_Sorter100|8308_  & \new_Sorter100|8309_ ;
  assign \new_Sorter100|8409_  = \new_Sorter100|8308_  | \new_Sorter100|8309_ ;
  assign \new_Sorter100|8410_  = \new_Sorter100|8310_  & \new_Sorter100|8311_ ;
  assign \new_Sorter100|8411_  = \new_Sorter100|8310_  | \new_Sorter100|8311_ ;
  assign \new_Sorter100|8412_  = \new_Sorter100|8312_  & \new_Sorter100|8313_ ;
  assign \new_Sorter100|8413_  = \new_Sorter100|8312_  | \new_Sorter100|8313_ ;
  assign \new_Sorter100|8414_  = \new_Sorter100|8314_  & \new_Sorter100|8315_ ;
  assign \new_Sorter100|8415_  = \new_Sorter100|8314_  | \new_Sorter100|8315_ ;
  assign \new_Sorter100|8416_  = \new_Sorter100|8316_  & \new_Sorter100|8317_ ;
  assign \new_Sorter100|8417_  = \new_Sorter100|8316_  | \new_Sorter100|8317_ ;
  assign \new_Sorter100|8418_  = \new_Sorter100|8318_  & \new_Sorter100|8319_ ;
  assign \new_Sorter100|8419_  = \new_Sorter100|8318_  | \new_Sorter100|8319_ ;
  assign \new_Sorter100|8420_  = \new_Sorter100|8320_  & \new_Sorter100|8321_ ;
  assign \new_Sorter100|8421_  = \new_Sorter100|8320_  | \new_Sorter100|8321_ ;
  assign \new_Sorter100|8422_  = \new_Sorter100|8322_  & \new_Sorter100|8323_ ;
  assign \new_Sorter100|8423_  = \new_Sorter100|8322_  | \new_Sorter100|8323_ ;
  assign \new_Sorter100|8424_  = \new_Sorter100|8324_  & \new_Sorter100|8325_ ;
  assign \new_Sorter100|8425_  = \new_Sorter100|8324_  | \new_Sorter100|8325_ ;
  assign \new_Sorter100|8426_  = \new_Sorter100|8326_  & \new_Sorter100|8327_ ;
  assign \new_Sorter100|8427_  = \new_Sorter100|8326_  | \new_Sorter100|8327_ ;
  assign \new_Sorter100|8428_  = \new_Sorter100|8328_  & \new_Sorter100|8329_ ;
  assign \new_Sorter100|8429_  = \new_Sorter100|8328_  | \new_Sorter100|8329_ ;
  assign \new_Sorter100|8430_  = \new_Sorter100|8330_  & \new_Sorter100|8331_ ;
  assign \new_Sorter100|8431_  = \new_Sorter100|8330_  | \new_Sorter100|8331_ ;
  assign \new_Sorter100|8432_  = \new_Sorter100|8332_  & \new_Sorter100|8333_ ;
  assign \new_Sorter100|8433_  = \new_Sorter100|8332_  | \new_Sorter100|8333_ ;
  assign \new_Sorter100|8434_  = \new_Sorter100|8334_  & \new_Sorter100|8335_ ;
  assign \new_Sorter100|8435_  = \new_Sorter100|8334_  | \new_Sorter100|8335_ ;
  assign \new_Sorter100|8436_  = \new_Sorter100|8336_  & \new_Sorter100|8337_ ;
  assign \new_Sorter100|8437_  = \new_Sorter100|8336_  | \new_Sorter100|8337_ ;
  assign \new_Sorter100|8438_  = \new_Sorter100|8338_  & \new_Sorter100|8339_ ;
  assign \new_Sorter100|8439_  = \new_Sorter100|8338_  | \new_Sorter100|8339_ ;
  assign \new_Sorter100|8440_  = \new_Sorter100|8340_  & \new_Sorter100|8341_ ;
  assign \new_Sorter100|8441_  = \new_Sorter100|8340_  | \new_Sorter100|8341_ ;
  assign \new_Sorter100|8442_  = \new_Sorter100|8342_  & \new_Sorter100|8343_ ;
  assign \new_Sorter100|8443_  = \new_Sorter100|8342_  | \new_Sorter100|8343_ ;
  assign \new_Sorter100|8444_  = \new_Sorter100|8344_  & \new_Sorter100|8345_ ;
  assign \new_Sorter100|8445_  = \new_Sorter100|8344_  | \new_Sorter100|8345_ ;
  assign \new_Sorter100|8446_  = \new_Sorter100|8346_  & \new_Sorter100|8347_ ;
  assign \new_Sorter100|8447_  = \new_Sorter100|8346_  | \new_Sorter100|8347_ ;
  assign \new_Sorter100|8448_  = \new_Sorter100|8348_  & \new_Sorter100|8349_ ;
  assign \new_Sorter100|8449_  = \new_Sorter100|8348_  | \new_Sorter100|8349_ ;
  assign \new_Sorter100|8450_  = \new_Sorter100|8350_  & \new_Sorter100|8351_ ;
  assign \new_Sorter100|8451_  = \new_Sorter100|8350_  | \new_Sorter100|8351_ ;
  assign \new_Sorter100|8452_  = \new_Sorter100|8352_  & \new_Sorter100|8353_ ;
  assign \new_Sorter100|8453_  = \new_Sorter100|8352_  | \new_Sorter100|8353_ ;
  assign \new_Sorter100|8454_  = \new_Sorter100|8354_  & \new_Sorter100|8355_ ;
  assign \new_Sorter100|8455_  = \new_Sorter100|8354_  | \new_Sorter100|8355_ ;
  assign \new_Sorter100|8456_  = \new_Sorter100|8356_  & \new_Sorter100|8357_ ;
  assign \new_Sorter100|8457_  = \new_Sorter100|8356_  | \new_Sorter100|8357_ ;
  assign \new_Sorter100|8458_  = \new_Sorter100|8358_  & \new_Sorter100|8359_ ;
  assign \new_Sorter100|8459_  = \new_Sorter100|8358_  | \new_Sorter100|8359_ ;
  assign \new_Sorter100|8460_  = \new_Sorter100|8360_  & \new_Sorter100|8361_ ;
  assign \new_Sorter100|8461_  = \new_Sorter100|8360_  | \new_Sorter100|8361_ ;
  assign \new_Sorter100|8462_  = \new_Sorter100|8362_  & \new_Sorter100|8363_ ;
  assign \new_Sorter100|8463_  = \new_Sorter100|8362_  | \new_Sorter100|8363_ ;
  assign \new_Sorter100|8464_  = \new_Sorter100|8364_  & \new_Sorter100|8365_ ;
  assign \new_Sorter100|8465_  = \new_Sorter100|8364_  | \new_Sorter100|8365_ ;
  assign \new_Sorter100|8466_  = \new_Sorter100|8366_  & \new_Sorter100|8367_ ;
  assign \new_Sorter100|8467_  = \new_Sorter100|8366_  | \new_Sorter100|8367_ ;
  assign \new_Sorter100|8468_  = \new_Sorter100|8368_  & \new_Sorter100|8369_ ;
  assign \new_Sorter100|8469_  = \new_Sorter100|8368_  | \new_Sorter100|8369_ ;
  assign \new_Sorter100|8470_  = \new_Sorter100|8370_  & \new_Sorter100|8371_ ;
  assign \new_Sorter100|8471_  = \new_Sorter100|8370_  | \new_Sorter100|8371_ ;
  assign \new_Sorter100|8472_  = \new_Sorter100|8372_  & \new_Sorter100|8373_ ;
  assign \new_Sorter100|8473_  = \new_Sorter100|8372_  | \new_Sorter100|8373_ ;
  assign \new_Sorter100|8474_  = \new_Sorter100|8374_  & \new_Sorter100|8375_ ;
  assign \new_Sorter100|8475_  = \new_Sorter100|8374_  | \new_Sorter100|8375_ ;
  assign \new_Sorter100|8476_  = \new_Sorter100|8376_  & \new_Sorter100|8377_ ;
  assign \new_Sorter100|8477_  = \new_Sorter100|8376_  | \new_Sorter100|8377_ ;
  assign \new_Sorter100|8478_  = \new_Sorter100|8378_  & \new_Sorter100|8379_ ;
  assign \new_Sorter100|8479_  = \new_Sorter100|8378_  | \new_Sorter100|8379_ ;
  assign \new_Sorter100|8480_  = \new_Sorter100|8380_  & \new_Sorter100|8381_ ;
  assign \new_Sorter100|8481_  = \new_Sorter100|8380_  | \new_Sorter100|8381_ ;
  assign \new_Sorter100|8482_  = \new_Sorter100|8382_  & \new_Sorter100|8383_ ;
  assign \new_Sorter100|8483_  = \new_Sorter100|8382_  | \new_Sorter100|8383_ ;
  assign \new_Sorter100|8484_  = \new_Sorter100|8384_  & \new_Sorter100|8385_ ;
  assign \new_Sorter100|8485_  = \new_Sorter100|8384_  | \new_Sorter100|8385_ ;
  assign \new_Sorter100|8486_  = \new_Sorter100|8386_  & \new_Sorter100|8387_ ;
  assign \new_Sorter100|8487_  = \new_Sorter100|8386_  | \new_Sorter100|8387_ ;
  assign \new_Sorter100|8488_  = \new_Sorter100|8388_  & \new_Sorter100|8389_ ;
  assign \new_Sorter100|8489_  = \new_Sorter100|8388_  | \new_Sorter100|8389_ ;
  assign \new_Sorter100|8490_  = \new_Sorter100|8390_  & \new_Sorter100|8391_ ;
  assign \new_Sorter100|8491_  = \new_Sorter100|8390_  | \new_Sorter100|8391_ ;
  assign \new_Sorter100|8492_  = \new_Sorter100|8392_  & \new_Sorter100|8393_ ;
  assign \new_Sorter100|8493_  = \new_Sorter100|8392_  | \new_Sorter100|8393_ ;
  assign \new_Sorter100|8494_  = \new_Sorter100|8394_  & \new_Sorter100|8395_ ;
  assign \new_Sorter100|8495_  = \new_Sorter100|8394_  | \new_Sorter100|8395_ ;
  assign \new_Sorter100|8496_  = \new_Sorter100|8396_  & \new_Sorter100|8397_ ;
  assign \new_Sorter100|8497_  = \new_Sorter100|8396_  | \new_Sorter100|8397_ ;
  assign \new_Sorter100|8498_  = \new_Sorter100|8398_  & \new_Sorter100|8399_ ;
  assign \new_Sorter100|8499_  = \new_Sorter100|8398_  | \new_Sorter100|8399_ ;
  assign \new_Sorter100|8500_  = \new_Sorter100|8400_ ;
  assign \new_Sorter100|8599_  = \new_Sorter100|8499_ ;
  assign \new_Sorter100|8501_  = \new_Sorter100|8401_  & \new_Sorter100|8402_ ;
  assign \new_Sorter100|8502_  = \new_Sorter100|8401_  | \new_Sorter100|8402_ ;
  assign \new_Sorter100|8503_  = \new_Sorter100|8403_  & \new_Sorter100|8404_ ;
  assign \new_Sorter100|8504_  = \new_Sorter100|8403_  | \new_Sorter100|8404_ ;
  assign \new_Sorter100|8505_  = \new_Sorter100|8405_  & \new_Sorter100|8406_ ;
  assign \new_Sorter100|8506_  = \new_Sorter100|8405_  | \new_Sorter100|8406_ ;
  assign \new_Sorter100|8507_  = \new_Sorter100|8407_  & \new_Sorter100|8408_ ;
  assign \new_Sorter100|8508_  = \new_Sorter100|8407_  | \new_Sorter100|8408_ ;
  assign \new_Sorter100|8509_  = \new_Sorter100|8409_  & \new_Sorter100|8410_ ;
  assign \new_Sorter100|8510_  = \new_Sorter100|8409_  | \new_Sorter100|8410_ ;
  assign \new_Sorter100|8511_  = \new_Sorter100|8411_  & \new_Sorter100|8412_ ;
  assign \new_Sorter100|8512_  = \new_Sorter100|8411_  | \new_Sorter100|8412_ ;
  assign \new_Sorter100|8513_  = \new_Sorter100|8413_  & \new_Sorter100|8414_ ;
  assign \new_Sorter100|8514_  = \new_Sorter100|8413_  | \new_Sorter100|8414_ ;
  assign \new_Sorter100|8515_  = \new_Sorter100|8415_  & \new_Sorter100|8416_ ;
  assign \new_Sorter100|8516_  = \new_Sorter100|8415_  | \new_Sorter100|8416_ ;
  assign \new_Sorter100|8517_  = \new_Sorter100|8417_  & \new_Sorter100|8418_ ;
  assign \new_Sorter100|8518_  = \new_Sorter100|8417_  | \new_Sorter100|8418_ ;
  assign \new_Sorter100|8519_  = \new_Sorter100|8419_  & \new_Sorter100|8420_ ;
  assign \new_Sorter100|8520_  = \new_Sorter100|8419_  | \new_Sorter100|8420_ ;
  assign \new_Sorter100|8521_  = \new_Sorter100|8421_  & \new_Sorter100|8422_ ;
  assign \new_Sorter100|8522_  = \new_Sorter100|8421_  | \new_Sorter100|8422_ ;
  assign \new_Sorter100|8523_  = \new_Sorter100|8423_  & \new_Sorter100|8424_ ;
  assign \new_Sorter100|8524_  = \new_Sorter100|8423_  | \new_Sorter100|8424_ ;
  assign \new_Sorter100|8525_  = \new_Sorter100|8425_  & \new_Sorter100|8426_ ;
  assign \new_Sorter100|8526_  = \new_Sorter100|8425_  | \new_Sorter100|8426_ ;
  assign \new_Sorter100|8527_  = \new_Sorter100|8427_  & \new_Sorter100|8428_ ;
  assign \new_Sorter100|8528_  = \new_Sorter100|8427_  | \new_Sorter100|8428_ ;
  assign \new_Sorter100|8529_  = \new_Sorter100|8429_  & \new_Sorter100|8430_ ;
  assign \new_Sorter100|8530_  = \new_Sorter100|8429_  | \new_Sorter100|8430_ ;
  assign \new_Sorter100|8531_  = \new_Sorter100|8431_  & \new_Sorter100|8432_ ;
  assign \new_Sorter100|8532_  = \new_Sorter100|8431_  | \new_Sorter100|8432_ ;
  assign \new_Sorter100|8533_  = \new_Sorter100|8433_  & \new_Sorter100|8434_ ;
  assign \new_Sorter100|8534_  = \new_Sorter100|8433_  | \new_Sorter100|8434_ ;
  assign \new_Sorter100|8535_  = \new_Sorter100|8435_  & \new_Sorter100|8436_ ;
  assign \new_Sorter100|8536_  = \new_Sorter100|8435_  | \new_Sorter100|8436_ ;
  assign \new_Sorter100|8537_  = \new_Sorter100|8437_  & \new_Sorter100|8438_ ;
  assign \new_Sorter100|8538_  = \new_Sorter100|8437_  | \new_Sorter100|8438_ ;
  assign \new_Sorter100|8539_  = \new_Sorter100|8439_  & \new_Sorter100|8440_ ;
  assign \new_Sorter100|8540_  = \new_Sorter100|8439_  | \new_Sorter100|8440_ ;
  assign \new_Sorter100|8541_  = \new_Sorter100|8441_  & \new_Sorter100|8442_ ;
  assign \new_Sorter100|8542_  = \new_Sorter100|8441_  | \new_Sorter100|8442_ ;
  assign \new_Sorter100|8543_  = \new_Sorter100|8443_  & \new_Sorter100|8444_ ;
  assign \new_Sorter100|8544_  = \new_Sorter100|8443_  | \new_Sorter100|8444_ ;
  assign \new_Sorter100|8545_  = \new_Sorter100|8445_  & \new_Sorter100|8446_ ;
  assign \new_Sorter100|8546_  = \new_Sorter100|8445_  | \new_Sorter100|8446_ ;
  assign \new_Sorter100|8547_  = \new_Sorter100|8447_  & \new_Sorter100|8448_ ;
  assign \new_Sorter100|8548_  = \new_Sorter100|8447_  | \new_Sorter100|8448_ ;
  assign \new_Sorter100|8549_  = \new_Sorter100|8449_  & \new_Sorter100|8450_ ;
  assign \new_Sorter100|8550_  = \new_Sorter100|8449_  | \new_Sorter100|8450_ ;
  assign \new_Sorter100|8551_  = \new_Sorter100|8451_  & \new_Sorter100|8452_ ;
  assign \new_Sorter100|8552_  = \new_Sorter100|8451_  | \new_Sorter100|8452_ ;
  assign \new_Sorter100|8553_  = \new_Sorter100|8453_  & \new_Sorter100|8454_ ;
  assign \new_Sorter100|8554_  = \new_Sorter100|8453_  | \new_Sorter100|8454_ ;
  assign \new_Sorter100|8555_  = \new_Sorter100|8455_  & \new_Sorter100|8456_ ;
  assign \new_Sorter100|8556_  = \new_Sorter100|8455_  | \new_Sorter100|8456_ ;
  assign \new_Sorter100|8557_  = \new_Sorter100|8457_  & \new_Sorter100|8458_ ;
  assign \new_Sorter100|8558_  = \new_Sorter100|8457_  | \new_Sorter100|8458_ ;
  assign \new_Sorter100|8559_  = \new_Sorter100|8459_  & \new_Sorter100|8460_ ;
  assign \new_Sorter100|8560_  = \new_Sorter100|8459_  | \new_Sorter100|8460_ ;
  assign \new_Sorter100|8561_  = \new_Sorter100|8461_  & \new_Sorter100|8462_ ;
  assign \new_Sorter100|8562_  = \new_Sorter100|8461_  | \new_Sorter100|8462_ ;
  assign \new_Sorter100|8563_  = \new_Sorter100|8463_  & \new_Sorter100|8464_ ;
  assign \new_Sorter100|8564_  = \new_Sorter100|8463_  | \new_Sorter100|8464_ ;
  assign \new_Sorter100|8565_  = \new_Sorter100|8465_  & \new_Sorter100|8466_ ;
  assign \new_Sorter100|8566_  = \new_Sorter100|8465_  | \new_Sorter100|8466_ ;
  assign \new_Sorter100|8567_  = \new_Sorter100|8467_  & \new_Sorter100|8468_ ;
  assign \new_Sorter100|8568_  = \new_Sorter100|8467_  | \new_Sorter100|8468_ ;
  assign \new_Sorter100|8569_  = \new_Sorter100|8469_  & \new_Sorter100|8470_ ;
  assign \new_Sorter100|8570_  = \new_Sorter100|8469_  | \new_Sorter100|8470_ ;
  assign \new_Sorter100|8571_  = \new_Sorter100|8471_  & \new_Sorter100|8472_ ;
  assign \new_Sorter100|8572_  = \new_Sorter100|8471_  | \new_Sorter100|8472_ ;
  assign \new_Sorter100|8573_  = \new_Sorter100|8473_  & \new_Sorter100|8474_ ;
  assign \new_Sorter100|8574_  = \new_Sorter100|8473_  | \new_Sorter100|8474_ ;
  assign \new_Sorter100|8575_  = \new_Sorter100|8475_  & \new_Sorter100|8476_ ;
  assign \new_Sorter100|8576_  = \new_Sorter100|8475_  | \new_Sorter100|8476_ ;
  assign \new_Sorter100|8577_  = \new_Sorter100|8477_  & \new_Sorter100|8478_ ;
  assign \new_Sorter100|8578_  = \new_Sorter100|8477_  | \new_Sorter100|8478_ ;
  assign \new_Sorter100|8579_  = \new_Sorter100|8479_  & \new_Sorter100|8480_ ;
  assign \new_Sorter100|8580_  = \new_Sorter100|8479_  | \new_Sorter100|8480_ ;
  assign \new_Sorter100|8581_  = \new_Sorter100|8481_  & \new_Sorter100|8482_ ;
  assign \new_Sorter100|8582_  = \new_Sorter100|8481_  | \new_Sorter100|8482_ ;
  assign \new_Sorter100|8583_  = \new_Sorter100|8483_  & \new_Sorter100|8484_ ;
  assign \new_Sorter100|8584_  = \new_Sorter100|8483_  | \new_Sorter100|8484_ ;
  assign \new_Sorter100|8585_  = \new_Sorter100|8485_  & \new_Sorter100|8486_ ;
  assign \new_Sorter100|8586_  = \new_Sorter100|8485_  | \new_Sorter100|8486_ ;
  assign \new_Sorter100|8587_  = \new_Sorter100|8487_  & \new_Sorter100|8488_ ;
  assign \new_Sorter100|8588_  = \new_Sorter100|8487_  | \new_Sorter100|8488_ ;
  assign \new_Sorter100|8589_  = \new_Sorter100|8489_  & \new_Sorter100|8490_ ;
  assign \new_Sorter100|8590_  = \new_Sorter100|8489_  | \new_Sorter100|8490_ ;
  assign \new_Sorter100|8591_  = \new_Sorter100|8491_  & \new_Sorter100|8492_ ;
  assign \new_Sorter100|8592_  = \new_Sorter100|8491_  | \new_Sorter100|8492_ ;
  assign \new_Sorter100|8593_  = \new_Sorter100|8493_  & \new_Sorter100|8494_ ;
  assign \new_Sorter100|8594_  = \new_Sorter100|8493_  | \new_Sorter100|8494_ ;
  assign \new_Sorter100|8595_  = \new_Sorter100|8495_  & \new_Sorter100|8496_ ;
  assign \new_Sorter100|8596_  = \new_Sorter100|8495_  | \new_Sorter100|8496_ ;
  assign \new_Sorter100|8597_  = \new_Sorter100|8497_  & \new_Sorter100|8498_ ;
  assign \new_Sorter100|8598_  = \new_Sorter100|8497_  | \new_Sorter100|8498_ ;
  assign \new_Sorter100|8600_  = \new_Sorter100|8500_  & \new_Sorter100|8501_ ;
  assign \new_Sorter100|8601_  = \new_Sorter100|8500_  | \new_Sorter100|8501_ ;
  assign \new_Sorter100|8602_  = \new_Sorter100|8502_  & \new_Sorter100|8503_ ;
  assign \new_Sorter100|8603_  = \new_Sorter100|8502_  | \new_Sorter100|8503_ ;
  assign \new_Sorter100|8604_  = \new_Sorter100|8504_  & \new_Sorter100|8505_ ;
  assign \new_Sorter100|8605_  = \new_Sorter100|8504_  | \new_Sorter100|8505_ ;
  assign \new_Sorter100|8606_  = \new_Sorter100|8506_  & \new_Sorter100|8507_ ;
  assign \new_Sorter100|8607_  = \new_Sorter100|8506_  | \new_Sorter100|8507_ ;
  assign \new_Sorter100|8608_  = \new_Sorter100|8508_  & \new_Sorter100|8509_ ;
  assign \new_Sorter100|8609_  = \new_Sorter100|8508_  | \new_Sorter100|8509_ ;
  assign \new_Sorter100|8610_  = \new_Sorter100|8510_  & \new_Sorter100|8511_ ;
  assign \new_Sorter100|8611_  = \new_Sorter100|8510_  | \new_Sorter100|8511_ ;
  assign \new_Sorter100|8612_  = \new_Sorter100|8512_  & \new_Sorter100|8513_ ;
  assign \new_Sorter100|8613_  = \new_Sorter100|8512_  | \new_Sorter100|8513_ ;
  assign \new_Sorter100|8614_  = \new_Sorter100|8514_  & \new_Sorter100|8515_ ;
  assign \new_Sorter100|8615_  = \new_Sorter100|8514_  | \new_Sorter100|8515_ ;
  assign \new_Sorter100|8616_  = \new_Sorter100|8516_  & \new_Sorter100|8517_ ;
  assign \new_Sorter100|8617_  = \new_Sorter100|8516_  | \new_Sorter100|8517_ ;
  assign \new_Sorter100|8618_  = \new_Sorter100|8518_  & \new_Sorter100|8519_ ;
  assign \new_Sorter100|8619_  = \new_Sorter100|8518_  | \new_Sorter100|8519_ ;
  assign \new_Sorter100|8620_  = \new_Sorter100|8520_  & \new_Sorter100|8521_ ;
  assign \new_Sorter100|8621_  = \new_Sorter100|8520_  | \new_Sorter100|8521_ ;
  assign \new_Sorter100|8622_  = \new_Sorter100|8522_  & \new_Sorter100|8523_ ;
  assign \new_Sorter100|8623_  = \new_Sorter100|8522_  | \new_Sorter100|8523_ ;
  assign \new_Sorter100|8624_  = \new_Sorter100|8524_  & \new_Sorter100|8525_ ;
  assign \new_Sorter100|8625_  = \new_Sorter100|8524_  | \new_Sorter100|8525_ ;
  assign \new_Sorter100|8626_  = \new_Sorter100|8526_  & \new_Sorter100|8527_ ;
  assign \new_Sorter100|8627_  = \new_Sorter100|8526_  | \new_Sorter100|8527_ ;
  assign \new_Sorter100|8628_  = \new_Sorter100|8528_  & \new_Sorter100|8529_ ;
  assign \new_Sorter100|8629_  = \new_Sorter100|8528_  | \new_Sorter100|8529_ ;
  assign \new_Sorter100|8630_  = \new_Sorter100|8530_  & \new_Sorter100|8531_ ;
  assign \new_Sorter100|8631_  = \new_Sorter100|8530_  | \new_Sorter100|8531_ ;
  assign \new_Sorter100|8632_  = \new_Sorter100|8532_  & \new_Sorter100|8533_ ;
  assign \new_Sorter100|8633_  = \new_Sorter100|8532_  | \new_Sorter100|8533_ ;
  assign \new_Sorter100|8634_  = \new_Sorter100|8534_  & \new_Sorter100|8535_ ;
  assign \new_Sorter100|8635_  = \new_Sorter100|8534_  | \new_Sorter100|8535_ ;
  assign \new_Sorter100|8636_  = \new_Sorter100|8536_  & \new_Sorter100|8537_ ;
  assign \new_Sorter100|8637_  = \new_Sorter100|8536_  | \new_Sorter100|8537_ ;
  assign \new_Sorter100|8638_  = \new_Sorter100|8538_  & \new_Sorter100|8539_ ;
  assign \new_Sorter100|8639_  = \new_Sorter100|8538_  | \new_Sorter100|8539_ ;
  assign \new_Sorter100|8640_  = \new_Sorter100|8540_  & \new_Sorter100|8541_ ;
  assign \new_Sorter100|8641_  = \new_Sorter100|8540_  | \new_Sorter100|8541_ ;
  assign \new_Sorter100|8642_  = \new_Sorter100|8542_  & \new_Sorter100|8543_ ;
  assign \new_Sorter100|8643_  = \new_Sorter100|8542_  | \new_Sorter100|8543_ ;
  assign \new_Sorter100|8644_  = \new_Sorter100|8544_  & \new_Sorter100|8545_ ;
  assign \new_Sorter100|8645_  = \new_Sorter100|8544_  | \new_Sorter100|8545_ ;
  assign \new_Sorter100|8646_  = \new_Sorter100|8546_  & \new_Sorter100|8547_ ;
  assign \new_Sorter100|8647_  = \new_Sorter100|8546_  | \new_Sorter100|8547_ ;
  assign \new_Sorter100|8648_  = \new_Sorter100|8548_  & \new_Sorter100|8549_ ;
  assign \new_Sorter100|8649_  = \new_Sorter100|8548_  | \new_Sorter100|8549_ ;
  assign \new_Sorter100|8650_  = \new_Sorter100|8550_  & \new_Sorter100|8551_ ;
  assign \new_Sorter100|8651_  = \new_Sorter100|8550_  | \new_Sorter100|8551_ ;
  assign \new_Sorter100|8652_  = \new_Sorter100|8552_  & \new_Sorter100|8553_ ;
  assign \new_Sorter100|8653_  = \new_Sorter100|8552_  | \new_Sorter100|8553_ ;
  assign \new_Sorter100|8654_  = \new_Sorter100|8554_  & \new_Sorter100|8555_ ;
  assign \new_Sorter100|8655_  = \new_Sorter100|8554_  | \new_Sorter100|8555_ ;
  assign \new_Sorter100|8656_  = \new_Sorter100|8556_  & \new_Sorter100|8557_ ;
  assign \new_Sorter100|8657_  = \new_Sorter100|8556_  | \new_Sorter100|8557_ ;
  assign \new_Sorter100|8658_  = \new_Sorter100|8558_  & \new_Sorter100|8559_ ;
  assign \new_Sorter100|8659_  = \new_Sorter100|8558_  | \new_Sorter100|8559_ ;
  assign \new_Sorter100|8660_  = \new_Sorter100|8560_  & \new_Sorter100|8561_ ;
  assign \new_Sorter100|8661_  = \new_Sorter100|8560_  | \new_Sorter100|8561_ ;
  assign \new_Sorter100|8662_  = \new_Sorter100|8562_  & \new_Sorter100|8563_ ;
  assign \new_Sorter100|8663_  = \new_Sorter100|8562_  | \new_Sorter100|8563_ ;
  assign \new_Sorter100|8664_  = \new_Sorter100|8564_  & \new_Sorter100|8565_ ;
  assign \new_Sorter100|8665_  = \new_Sorter100|8564_  | \new_Sorter100|8565_ ;
  assign \new_Sorter100|8666_  = \new_Sorter100|8566_  & \new_Sorter100|8567_ ;
  assign \new_Sorter100|8667_  = \new_Sorter100|8566_  | \new_Sorter100|8567_ ;
  assign \new_Sorter100|8668_  = \new_Sorter100|8568_  & \new_Sorter100|8569_ ;
  assign \new_Sorter100|8669_  = \new_Sorter100|8568_  | \new_Sorter100|8569_ ;
  assign \new_Sorter100|8670_  = \new_Sorter100|8570_  & \new_Sorter100|8571_ ;
  assign \new_Sorter100|8671_  = \new_Sorter100|8570_  | \new_Sorter100|8571_ ;
  assign \new_Sorter100|8672_  = \new_Sorter100|8572_  & \new_Sorter100|8573_ ;
  assign \new_Sorter100|8673_  = \new_Sorter100|8572_  | \new_Sorter100|8573_ ;
  assign \new_Sorter100|8674_  = \new_Sorter100|8574_  & \new_Sorter100|8575_ ;
  assign \new_Sorter100|8675_  = \new_Sorter100|8574_  | \new_Sorter100|8575_ ;
  assign \new_Sorter100|8676_  = \new_Sorter100|8576_  & \new_Sorter100|8577_ ;
  assign \new_Sorter100|8677_  = \new_Sorter100|8576_  | \new_Sorter100|8577_ ;
  assign \new_Sorter100|8678_  = \new_Sorter100|8578_  & \new_Sorter100|8579_ ;
  assign \new_Sorter100|8679_  = \new_Sorter100|8578_  | \new_Sorter100|8579_ ;
  assign \new_Sorter100|8680_  = \new_Sorter100|8580_  & \new_Sorter100|8581_ ;
  assign \new_Sorter100|8681_  = \new_Sorter100|8580_  | \new_Sorter100|8581_ ;
  assign \new_Sorter100|8682_  = \new_Sorter100|8582_  & \new_Sorter100|8583_ ;
  assign \new_Sorter100|8683_  = \new_Sorter100|8582_  | \new_Sorter100|8583_ ;
  assign \new_Sorter100|8684_  = \new_Sorter100|8584_  & \new_Sorter100|8585_ ;
  assign \new_Sorter100|8685_  = \new_Sorter100|8584_  | \new_Sorter100|8585_ ;
  assign \new_Sorter100|8686_  = \new_Sorter100|8586_  & \new_Sorter100|8587_ ;
  assign \new_Sorter100|8687_  = \new_Sorter100|8586_  | \new_Sorter100|8587_ ;
  assign \new_Sorter100|8688_  = \new_Sorter100|8588_  & \new_Sorter100|8589_ ;
  assign \new_Sorter100|8689_  = \new_Sorter100|8588_  | \new_Sorter100|8589_ ;
  assign \new_Sorter100|8690_  = \new_Sorter100|8590_  & \new_Sorter100|8591_ ;
  assign \new_Sorter100|8691_  = \new_Sorter100|8590_  | \new_Sorter100|8591_ ;
  assign \new_Sorter100|8692_  = \new_Sorter100|8592_  & \new_Sorter100|8593_ ;
  assign \new_Sorter100|8693_  = \new_Sorter100|8592_  | \new_Sorter100|8593_ ;
  assign \new_Sorter100|8694_  = \new_Sorter100|8594_  & \new_Sorter100|8595_ ;
  assign \new_Sorter100|8695_  = \new_Sorter100|8594_  | \new_Sorter100|8595_ ;
  assign \new_Sorter100|8696_  = \new_Sorter100|8596_  & \new_Sorter100|8597_ ;
  assign \new_Sorter100|8697_  = \new_Sorter100|8596_  | \new_Sorter100|8597_ ;
  assign \new_Sorter100|8698_  = \new_Sorter100|8598_  & \new_Sorter100|8599_ ;
  assign \new_Sorter100|8699_  = \new_Sorter100|8598_  | \new_Sorter100|8599_ ;
  assign \new_Sorter100|8700_  = \new_Sorter100|8600_ ;
  assign \new_Sorter100|8799_  = \new_Sorter100|8699_ ;
  assign \new_Sorter100|8701_  = \new_Sorter100|8601_  & \new_Sorter100|8602_ ;
  assign \new_Sorter100|8702_  = \new_Sorter100|8601_  | \new_Sorter100|8602_ ;
  assign \new_Sorter100|8703_  = \new_Sorter100|8603_  & \new_Sorter100|8604_ ;
  assign \new_Sorter100|8704_  = \new_Sorter100|8603_  | \new_Sorter100|8604_ ;
  assign \new_Sorter100|8705_  = \new_Sorter100|8605_  & \new_Sorter100|8606_ ;
  assign \new_Sorter100|8706_  = \new_Sorter100|8605_  | \new_Sorter100|8606_ ;
  assign \new_Sorter100|8707_  = \new_Sorter100|8607_  & \new_Sorter100|8608_ ;
  assign \new_Sorter100|8708_  = \new_Sorter100|8607_  | \new_Sorter100|8608_ ;
  assign \new_Sorter100|8709_  = \new_Sorter100|8609_  & \new_Sorter100|8610_ ;
  assign \new_Sorter100|8710_  = \new_Sorter100|8609_  | \new_Sorter100|8610_ ;
  assign \new_Sorter100|8711_  = \new_Sorter100|8611_  & \new_Sorter100|8612_ ;
  assign \new_Sorter100|8712_  = \new_Sorter100|8611_  | \new_Sorter100|8612_ ;
  assign \new_Sorter100|8713_  = \new_Sorter100|8613_  & \new_Sorter100|8614_ ;
  assign \new_Sorter100|8714_  = \new_Sorter100|8613_  | \new_Sorter100|8614_ ;
  assign \new_Sorter100|8715_  = \new_Sorter100|8615_  & \new_Sorter100|8616_ ;
  assign \new_Sorter100|8716_  = \new_Sorter100|8615_  | \new_Sorter100|8616_ ;
  assign \new_Sorter100|8717_  = \new_Sorter100|8617_  & \new_Sorter100|8618_ ;
  assign \new_Sorter100|8718_  = \new_Sorter100|8617_  | \new_Sorter100|8618_ ;
  assign \new_Sorter100|8719_  = \new_Sorter100|8619_  & \new_Sorter100|8620_ ;
  assign \new_Sorter100|8720_  = \new_Sorter100|8619_  | \new_Sorter100|8620_ ;
  assign \new_Sorter100|8721_  = \new_Sorter100|8621_  & \new_Sorter100|8622_ ;
  assign \new_Sorter100|8722_  = \new_Sorter100|8621_  | \new_Sorter100|8622_ ;
  assign \new_Sorter100|8723_  = \new_Sorter100|8623_  & \new_Sorter100|8624_ ;
  assign \new_Sorter100|8724_  = \new_Sorter100|8623_  | \new_Sorter100|8624_ ;
  assign \new_Sorter100|8725_  = \new_Sorter100|8625_  & \new_Sorter100|8626_ ;
  assign \new_Sorter100|8726_  = \new_Sorter100|8625_  | \new_Sorter100|8626_ ;
  assign \new_Sorter100|8727_  = \new_Sorter100|8627_  & \new_Sorter100|8628_ ;
  assign \new_Sorter100|8728_  = \new_Sorter100|8627_  | \new_Sorter100|8628_ ;
  assign \new_Sorter100|8729_  = \new_Sorter100|8629_  & \new_Sorter100|8630_ ;
  assign \new_Sorter100|8730_  = \new_Sorter100|8629_  | \new_Sorter100|8630_ ;
  assign \new_Sorter100|8731_  = \new_Sorter100|8631_  & \new_Sorter100|8632_ ;
  assign \new_Sorter100|8732_  = \new_Sorter100|8631_  | \new_Sorter100|8632_ ;
  assign \new_Sorter100|8733_  = \new_Sorter100|8633_  & \new_Sorter100|8634_ ;
  assign \new_Sorter100|8734_  = \new_Sorter100|8633_  | \new_Sorter100|8634_ ;
  assign \new_Sorter100|8735_  = \new_Sorter100|8635_  & \new_Sorter100|8636_ ;
  assign \new_Sorter100|8736_  = \new_Sorter100|8635_  | \new_Sorter100|8636_ ;
  assign \new_Sorter100|8737_  = \new_Sorter100|8637_  & \new_Sorter100|8638_ ;
  assign \new_Sorter100|8738_  = \new_Sorter100|8637_  | \new_Sorter100|8638_ ;
  assign \new_Sorter100|8739_  = \new_Sorter100|8639_  & \new_Sorter100|8640_ ;
  assign \new_Sorter100|8740_  = \new_Sorter100|8639_  | \new_Sorter100|8640_ ;
  assign \new_Sorter100|8741_  = \new_Sorter100|8641_  & \new_Sorter100|8642_ ;
  assign \new_Sorter100|8742_  = \new_Sorter100|8641_  | \new_Sorter100|8642_ ;
  assign \new_Sorter100|8743_  = \new_Sorter100|8643_  & \new_Sorter100|8644_ ;
  assign \new_Sorter100|8744_  = \new_Sorter100|8643_  | \new_Sorter100|8644_ ;
  assign \new_Sorter100|8745_  = \new_Sorter100|8645_  & \new_Sorter100|8646_ ;
  assign \new_Sorter100|8746_  = \new_Sorter100|8645_  | \new_Sorter100|8646_ ;
  assign \new_Sorter100|8747_  = \new_Sorter100|8647_  & \new_Sorter100|8648_ ;
  assign \new_Sorter100|8748_  = \new_Sorter100|8647_  | \new_Sorter100|8648_ ;
  assign \new_Sorter100|8749_  = \new_Sorter100|8649_  & \new_Sorter100|8650_ ;
  assign \new_Sorter100|8750_  = \new_Sorter100|8649_  | \new_Sorter100|8650_ ;
  assign \new_Sorter100|8751_  = \new_Sorter100|8651_  & \new_Sorter100|8652_ ;
  assign \new_Sorter100|8752_  = \new_Sorter100|8651_  | \new_Sorter100|8652_ ;
  assign \new_Sorter100|8753_  = \new_Sorter100|8653_  & \new_Sorter100|8654_ ;
  assign \new_Sorter100|8754_  = \new_Sorter100|8653_  | \new_Sorter100|8654_ ;
  assign \new_Sorter100|8755_  = \new_Sorter100|8655_  & \new_Sorter100|8656_ ;
  assign \new_Sorter100|8756_  = \new_Sorter100|8655_  | \new_Sorter100|8656_ ;
  assign \new_Sorter100|8757_  = \new_Sorter100|8657_  & \new_Sorter100|8658_ ;
  assign \new_Sorter100|8758_  = \new_Sorter100|8657_  | \new_Sorter100|8658_ ;
  assign \new_Sorter100|8759_  = \new_Sorter100|8659_  & \new_Sorter100|8660_ ;
  assign \new_Sorter100|8760_  = \new_Sorter100|8659_  | \new_Sorter100|8660_ ;
  assign \new_Sorter100|8761_  = \new_Sorter100|8661_  & \new_Sorter100|8662_ ;
  assign \new_Sorter100|8762_  = \new_Sorter100|8661_  | \new_Sorter100|8662_ ;
  assign \new_Sorter100|8763_  = \new_Sorter100|8663_  & \new_Sorter100|8664_ ;
  assign \new_Sorter100|8764_  = \new_Sorter100|8663_  | \new_Sorter100|8664_ ;
  assign \new_Sorter100|8765_  = \new_Sorter100|8665_  & \new_Sorter100|8666_ ;
  assign \new_Sorter100|8766_  = \new_Sorter100|8665_  | \new_Sorter100|8666_ ;
  assign \new_Sorter100|8767_  = \new_Sorter100|8667_  & \new_Sorter100|8668_ ;
  assign \new_Sorter100|8768_  = \new_Sorter100|8667_  | \new_Sorter100|8668_ ;
  assign \new_Sorter100|8769_  = \new_Sorter100|8669_  & \new_Sorter100|8670_ ;
  assign \new_Sorter100|8770_  = \new_Sorter100|8669_  | \new_Sorter100|8670_ ;
  assign \new_Sorter100|8771_  = \new_Sorter100|8671_  & \new_Sorter100|8672_ ;
  assign \new_Sorter100|8772_  = \new_Sorter100|8671_  | \new_Sorter100|8672_ ;
  assign \new_Sorter100|8773_  = \new_Sorter100|8673_  & \new_Sorter100|8674_ ;
  assign \new_Sorter100|8774_  = \new_Sorter100|8673_  | \new_Sorter100|8674_ ;
  assign \new_Sorter100|8775_  = \new_Sorter100|8675_  & \new_Sorter100|8676_ ;
  assign \new_Sorter100|8776_  = \new_Sorter100|8675_  | \new_Sorter100|8676_ ;
  assign \new_Sorter100|8777_  = \new_Sorter100|8677_  & \new_Sorter100|8678_ ;
  assign \new_Sorter100|8778_  = \new_Sorter100|8677_  | \new_Sorter100|8678_ ;
  assign \new_Sorter100|8779_  = \new_Sorter100|8679_  & \new_Sorter100|8680_ ;
  assign \new_Sorter100|8780_  = \new_Sorter100|8679_  | \new_Sorter100|8680_ ;
  assign \new_Sorter100|8781_  = \new_Sorter100|8681_  & \new_Sorter100|8682_ ;
  assign \new_Sorter100|8782_  = \new_Sorter100|8681_  | \new_Sorter100|8682_ ;
  assign \new_Sorter100|8783_  = \new_Sorter100|8683_  & \new_Sorter100|8684_ ;
  assign \new_Sorter100|8784_  = \new_Sorter100|8683_  | \new_Sorter100|8684_ ;
  assign \new_Sorter100|8785_  = \new_Sorter100|8685_  & \new_Sorter100|8686_ ;
  assign \new_Sorter100|8786_  = \new_Sorter100|8685_  | \new_Sorter100|8686_ ;
  assign \new_Sorter100|8787_  = \new_Sorter100|8687_  & \new_Sorter100|8688_ ;
  assign \new_Sorter100|8788_  = \new_Sorter100|8687_  | \new_Sorter100|8688_ ;
  assign \new_Sorter100|8789_  = \new_Sorter100|8689_  & \new_Sorter100|8690_ ;
  assign \new_Sorter100|8790_  = \new_Sorter100|8689_  | \new_Sorter100|8690_ ;
  assign \new_Sorter100|8791_  = \new_Sorter100|8691_  & \new_Sorter100|8692_ ;
  assign \new_Sorter100|8792_  = \new_Sorter100|8691_  | \new_Sorter100|8692_ ;
  assign \new_Sorter100|8793_  = \new_Sorter100|8693_  & \new_Sorter100|8694_ ;
  assign \new_Sorter100|8794_  = \new_Sorter100|8693_  | \new_Sorter100|8694_ ;
  assign \new_Sorter100|8795_  = \new_Sorter100|8695_  & \new_Sorter100|8696_ ;
  assign \new_Sorter100|8796_  = \new_Sorter100|8695_  | \new_Sorter100|8696_ ;
  assign \new_Sorter100|8797_  = \new_Sorter100|8697_  & \new_Sorter100|8698_ ;
  assign \new_Sorter100|8798_  = \new_Sorter100|8697_  | \new_Sorter100|8698_ ;
  assign \new_Sorter100|8800_  = \new_Sorter100|8700_  & \new_Sorter100|8701_ ;
  assign \new_Sorter100|8801_  = \new_Sorter100|8700_  | \new_Sorter100|8701_ ;
  assign \new_Sorter100|8802_  = \new_Sorter100|8702_  & \new_Sorter100|8703_ ;
  assign \new_Sorter100|8803_  = \new_Sorter100|8702_  | \new_Sorter100|8703_ ;
  assign \new_Sorter100|8804_  = \new_Sorter100|8704_  & \new_Sorter100|8705_ ;
  assign \new_Sorter100|8805_  = \new_Sorter100|8704_  | \new_Sorter100|8705_ ;
  assign \new_Sorter100|8806_  = \new_Sorter100|8706_  & \new_Sorter100|8707_ ;
  assign \new_Sorter100|8807_  = \new_Sorter100|8706_  | \new_Sorter100|8707_ ;
  assign \new_Sorter100|8808_  = \new_Sorter100|8708_  & \new_Sorter100|8709_ ;
  assign \new_Sorter100|8809_  = \new_Sorter100|8708_  | \new_Sorter100|8709_ ;
  assign \new_Sorter100|8810_  = \new_Sorter100|8710_  & \new_Sorter100|8711_ ;
  assign \new_Sorter100|8811_  = \new_Sorter100|8710_  | \new_Sorter100|8711_ ;
  assign \new_Sorter100|8812_  = \new_Sorter100|8712_  & \new_Sorter100|8713_ ;
  assign \new_Sorter100|8813_  = \new_Sorter100|8712_  | \new_Sorter100|8713_ ;
  assign \new_Sorter100|8814_  = \new_Sorter100|8714_  & \new_Sorter100|8715_ ;
  assign \new_Sorter100|8815_  = \new_Sorter100|8714_  | \new_Sorter100|8715_ ;
  assign \new_Sorter100|8816_  = \new_Sorter100|8716_  & \new_Sorter100|8717_ ;
  assign \new_Sorter100|8817_  = \new_Sorter100|8716_  | \new_Sorter100|8717_ ;
  assign \new_Sorter100|8818_  = \new_Sorter100|8718_  & \new_Sorter100|8719_ ;
  assign \new_Sorter100|8819_  = \new_Sorter100|8718_  | \new_Sorter100|8719_ ;
  assign \new_Sorter100|8820_  = \new_Sorter100|8720_  & \new_Sorter100|8721_ ;
  assign \new_Sorter100|8821_  = \new_Sorter100|8720_  | \new_Sorter100|8721_ ;
  assign \new_Sorter100|8822_  = \new_Sorter100|8722_  & \new_Sorter100|8723_ ;
  assign \new_Sorter100|8823_  = \new_Sorter100|8722_  | \new_Sorter100|8723_ ;
  assign \new_Sorter100|8824_  = \new_Sorter100|8724_  & \new_Sorter100|8725_ ;
  assign \new_Sorter100|8825_  = \new_Sorter100|8724_  | \new_Sorter100|8725_ ;
  assign \new_Sorter100|8826_  = \new_Sorter100|8726_  & \new_Sorter100|8727_ ;
  assign \new_Sorter100|8827_  = \new_Sorter100|8726_  | \new_Sorter100|8727_ ;
  assign \new_Sorter100|8828_  = \new_Sorter100|8728_  & \new_Sorter100|8729_ ;
  assign \new_Sorter100|8829_  = \new_Sorter100|8728_  | \new_Sorter100|8729_ ;
  assign \new_Sorter100|8830_  = \new_Sorter100|8730_  & \new_Sorter100|8731_ ;
  assign \new_Sorter100|8831_  = \new_Sorter100|8730_  | \new_Sorter100|8731_ ;
  assign \new_Sorter100|8832_  = \new_Sorter100|8732_  & \new_Sorter100|8733_ ;
  assign \new_Sorter100|8833_  = \new_Sorter100|8732_  | \new_Sorter100|8733_ ;
  assign \new_Sorter100|8834_  = \new_Sorter100|8734_  & \new_Sorter100|8735_ ;
  assign \new_Sorter100|8835_  = \new_Sorter100|8734_  | \new_Sorter100|8735_ ;
  assign \new_Sorter100|8836_  = \new_Sorter100|8736_  & \new_Sorter100|8737_ ;
  assign \new_Sorter100|8837_  = \new_Sorter100|8736_  | \new_Sorter100|8737_ ;
  assign \new_Sorter100|8838_  = \new_Sorter100|8738_  & \new_Sorter100|8739_ ;
  assign \new_Sorter100|8839_  = \new_Sorter100|8738_  | \new_Sorter100|8739_ ;
  assign \new_Sorter100|8840_  = \new_Sorter100|8740_  & \new_Sorter100|8741_ ;
  assign \new_Sorter100|8841_  = \new_Sorter100|8740_  | \new_Sorter100|8741_ ;
  assign \new_Sorter100|8842_  = \new_Sorter100|8742_  & \new_Sorter100|8743_ ;
  assign \new_Sorter100|8843_  = \new_Sorter100|8742_  | \new_Sorter100|8743_ ;
  assign \new_Sorter100|8844_  = \new_Sorter100|8744_  & \new_Sorter100|8745_ ;
  assign \new_Sorter100|8845_  = \new_Sorter100|8744_  | \new_Sorter100|8745_ ;
  assign \new_Sorter100|8846_  = \new_Sorter100|8746_  & \new_Sorter100|8747_ ;
  assign \new_Sorter100|8847_  = \new_Sorter100|8746_  | \new_Sorter100|8747_ ;
  assign \new_Sorter100|8848_  = \new_Sorter100|8748_  & \new_Sorter100|8749_ ;
  assign \new_Sorter100|8849_  = \new_Sorter100|8748_  | \new_Sorter100|8749_ ;
  assign \new_Sorter100|8850_  = \new_Sorter100|8750_  & \new_Sorter100|8751_ ;
  assign \new_Sorter100|8851_  = \new_Sorter100|8750_  | \new_Sorter100|8751_ ;
  assign \new_Sorter100|8852_  = \new_Sorter100|8752_  & \new_Sorter100|8753_ ;
  assign \new_Sorter100|8853_  = \new_Sorter100|8752_  | \new_Sorter100|8753_ ;
  assign \new_Sorter100|8854_  = \new_Sorter100|8754_  & \new_Sorter100|8755_ ;
  assign \new_Sorter100|8855_  = \new_Sorter100|8754_  | \new_Sorter100|8755_ ;
  assign \new_Sorter100|8856_  = \new_Sorter100|8756_  & \new_Sorter100|8757_ ;
  assign \new_Sorter100|8857_  = \new_Sorter100|8756_  | \new_Sorter100|8757_ ;
  assign \new_Sorter100|8858_  = \new_Sorter100|8758_  & \new_Sorter100|8759_ ;
  assign \new_Sorter100|8859_  = \new_Sorter100|8758_  | \new_Sorter100|8759_ ;
  assign \new_Sorter100|8860_  = \new_Sorter100|8760_  & \new_Sorter100|8761_ ;
  assign \new_Sorter100|8861_  = \new_Sorter100|8760_  | \new_Sorter100|8761_ ;
  assign \new_Sorter100|8862_  = \new_Sorter100|8762_  & \new_Sorter100|8763_ ;
  assign \new_Sorter100|8863_  = \new_Sorter100|8762_  | \new_Sorter100|8763_ ;
  assign \new_Sorter100|8864_  = \new_Sorter100|8764_  & \new_Sorter100|8765_ ;
  assign \new_Sorter100|8865_  = \new_Sorter100|8764_  | \new_Sorter100|8765_ ;
  assign \new_Sorter100|8866_  = \new_Sorter100|8766_  & \new_Sorter100|8767_ ;
  assign \new_Sorter100|8867_  = \new_Sorter100|8766_  | \new_Sorter100|8767_ ;
  assign \new_Sorter100|8868_  = \new_Sorter100|8768_  & \new_Sorter100|8769_ ;
  assign \new_Sorter100|8869_  = \new_Sorter100|8768_  | \new_Sorter100|8769_ ;
  assign \new_Sorter100|8870_  = \new_Sorter100|8770_  & \new_Sorter100|8771_ ;
  assign \new_Sorter100|8871_  = \new_Sorter100|8770_  | \new_Sorter100|8771_ ;
  assign \new_Sorter100|8872_  = \new_Sorter100|8772_  & \new_Sorter100|8773_ ;
  assign \new_Sorter100|8873_  = \new_Sorter100|8772_  | \new_Sorter100|8773_ ;
  assign \new_Sorter100|8874_  = \new_Sorter100|8774_  & \new_Sorter100|8775_ ;
  assign \new_Sorter100|8875_  = \new_Sorter100|8774_  | \new_Sorter100|8775_ ;
  assign \new_Sorter100|8876_  = \new_Sorter100|8776_  & \new_Sorter100|8777_ ;
  assign \new_Sorter100|8877_  = \new_Sorter100|8776_  | \new_Sorter100|8777_ ;
  assign \new_Sorter100|8878_  = \new_Sorter100|8778_  & \new_Sorter100|8779_ ;
  assign \new_Sorter100|8879_  = \new_Sorter100|8778_  | \new_Sorter100|8779_ ;
  assign \new_Sorter100|8880_  = \new_Sorter100|8780_  & \new_Sorter100|8781_ ;
  assign \new_Sorter100|8881_  = \new_Sorter100|8780_  | \new_Sorter100|8781_ ;
  assign \new_Sorter100|8882_  = \new_Sorter100|8782_  & \new_Sorter100|8783_ ;
  assign \new_Sorter100|8883_  = \new_Sorter100|8782_  | \new_Sorter100|8783_ ;
  assign \new_Sorter100|8884_  = \new_Sorter100|8784_  & \new_Sorter100|8785_ ;
  assign \new_Sorter100|8885_  = \new_Sorter100|8784_  | \new_Sorter100|8785_ ;
  assign \new_Sorter100|8886_  = \new_Sorter100|8786_  & \new_Sorter100|8787_ ;
  assign \new_Sorter100|8887_  = \new_Sorter100|8786_  | \new_Sorter100|8787_ ;
  assign \new_Sorter100|8888_  = \new_Sorter100|8788_  & \new_Sorter100|8789_ ;
  assign \new_Sorter100|8889_  = \new_Sorter100|8788_  | \new_Sorter100|8789_ ;
  assign \new_Sorter100|8890_  = \new_Sorter100|8790_  & \new_Sorter100|8791_ ;
  assign \new_Sorter100|8891_  = \new_Sorter100|8790_  | \new_Sorter100|8791_ ;
  assign \new_Sorter100|8892_  = \new_Sorter100|8792_  & \new_Sorter100|8793_ ;
  assign \new_Sorter100|8893_  = \new_Sorter100|8792_  | \new_Sorter100|8793_ ;
  assign \new_Sorter100|8894_  = \new_Sorter100|8794_  & \new_Sorter100|8795_ ;
  assign \new_Sorter100|8895_  = \new_Sorter100|8794_  | \new_Sorter100|8795_ ;
  assign \new_Sorter100|8896_  = \new_Sorter100|8796_  & \new_Sorter100|8797_ ;
  assign \new_Sorter100|8897_  = \new_Sorter100|8796_  | \new_Sorter100|8797_ ;
  assign \new_Sorter100|8898_  = \new_Sorter100|8798_  & \new_Sorter100|8799_ ;
  assign \new_Sorter100|8899_  = \new_Sorter100|8798_  | \new_Sorter100|8799_ ;
  assign \new_Sorter100|8900_  = \new_Sorter100|8800_ ;
  assign \new_Sorter100|8999_  = \new_Sorter100|8899_ ;
  assign \new_Sorter100|8901_  = \new_Sorter100|8801_  & \new_Sorter100|8802_ ;
  assign \new_Sorter100|8902_  = \new_Sorter100|8801_  | \new_Sorter100|8802_ ;
  assign \new_Sorter100|8903_  = \new_Sorter100|8803_  & \new_Sorter100|8804_ ;
  assign \new_Sorter100|8904_  = \new_Sorter100|8803_  | \new_Sorter100|8804_ ;
  assign \new_Sorter100|8905_  = \new_Sorter100|8805_  & \new_Sorter100|8806_ ;
  assign \new_Sorter100|8906_  = \new_Sorter100|8805_  | \new_Sorter100|8806_ ;
  assign \new_Sorter100|8907_  = \new_Sorter100|8807_  & \new_Sorter100|8808_ ;
  assign \new_Sorter100|8908_  = \new_Sorter100|8807_  | \new_Sorter100|8808_ ;
  assign \new_Sorter100|8909_  = \new_Sorter100|8809_  & \new_Sorter100|8810_ ;
  assign \new_Sorter100|8910_  = \new_Sorter100|8809_  | \new_Sorter100|8810_ ;
  assign \new_Sorter100|8911_  = \new_Sorter100|8811_  & \new_Sorter100|8812_ ;
  assign \new_Sorter100|8912_  = \new_Sorter100|8811_  | \new_Sorter100|8812_ ;
  assign \new_Sorter100|8913_  = \new_Sorter100|8813_  & \new_Sorter100|8814_ ;
  assign \new_Sorter100|8914_  = \new_Sorter100|8813_  | \new_Sorter100|8814_ ;
  assign \new_Sorter100|8915_  = \new_Sorter100|8815_  & \new_Sorter100|8816_ ;
  assign \new_Sorter100|8916_  = \new_Sorter100|8815_  | \new_Sorter100|8816_ ;
  assign \new_Sorter100|8917_  = \new_Sorter100|8817_  & \new_Sorter100|8818_ ;
  assign \new_Sorter100|8918_  = \new_Sorter100|8817_  | \new_Sorter100|8818_ ;
  assign \new_Sorter100|8919_  = \new_Sorter100|8819_  & \new_Sorter100|8820_ ;
  assign \new_Sorter100|8920_  = \new_Sorter100|8819_  | \new_Sorter100|8820_ ;
  assign \new_Sorter100|8921_  = \new_Sorter100|8821_  & \new_Sorter100|8822_ ;
  assign \new_Sorter100|8922_  = \new_Sorter100|8821_  | \new_Sorter100|8822_ ;
  assign \new_Sorter100|8923_  = \new_Sorter100|8823_  & \new_Sorter100|8824_ ;
  assign \new_Sorter100|8924_  = \new_Sorter100|8823_  | \new_Sorter100|8824_ ;
  assign \new_Sorter100|8925_  = \new_Sorter100|8825_  & \new_Sorter100|8826_ ;
  assign \new_Sorter100|8926_  = \new_Sorter100|8825_  | \new_Sorter100|8826_ ;
  assign \new_Sorter100|8927_  = \new_Sorter100|8827_  & \new_Sorter100|8828_ ;
  assign \new_Sorter100|8928_  = \new_Sorter100|8827_  | \new_Sorter100|8828_ ;
  assign \new_Sorter100|8929_  = \new_Sorter100|8829_  & \new_Sorter100|8830_ ;
  assign \new_Sorter100|8930_  = \new_Sorter100|8829_  | \new_Sorter100|8830_ ;
  assign \new_Sorter100|8931_  = \new_Sorter100|8831_  & \new_Sorter100|8832_ ;
  assign \new_Sorter100|8932_  = \new_Sorter100|8831_  | \new_Sorter100|8832_ ;
  assign \new_Sorter100|8933_  = \new_Sorter100|8833_  & \new_Sorter100|8834_ ;
  assign \new_Sorter100|8934_  = \new_Sorter100|8833_  | \new_Sorter100|8834_ ;
  assign \new_Sorter100|8935_  = \new_Sorter100|8835_  & \new_Sorter100|8836_ ;
  assign \new_Sorter100|8936_  = \new_Sorter100|8835_  | \new_Sorter100|8836_ ;
  assign \new_Sorter100|8937_  = \new_Sorter100|8837_  & \new_Sorter100|8838_ ;
  assign \new_Sorter100|8938_  = \new_Sorter100|8837_  | \new_Sorter100|8838_ ;
  assign \new_Sorter100|8939_  = \new_Sorter100|8839_  & \new_Sorter100|8840_ ;
  assign \new_Sorter100|8940_  = \new_Sorter100|8839_  | \new_Sorter100|8840_ ;
  assign \new_Sorter100|8941_  = \new_Sorter100|8841_  & \new_Sorter100|8842_ ;
  assign \new_Sorter100|8942_  = \new_Sorter100|8841_  | \new_Sorter100|8842_ ;
  assign \new_Sorter100|8943_  = \new_Sorter100|8843_  & \new_Sorter100|8844_ ;
  assign \new_Sorter100|8944_  = \new_Sorter100|8843_  | \new_Sorter100|8844_ ;
  assign \new_Sorter100|8945_  = \new_Sorter100|8845_  & \new_Sorter100|8846_ ;
  assign \new_Sorter100|8946_  = \new_Sorter100|8845_  | \new_Sorter100|8846_ ;
  assign \new_Sorter100|8947_  = \new_Sorter100|8847_  & \new_Sorter100|8848_ ;
  assign \new_Sorter100|8948_  = \new_Sorter100|8847_  | \new_Sorter100|8848_ ;
  assign \new_Sorter100|8949_  = \new_Sorter100|8849_  & \new_Sorter100|8850_ ;
  assign \new_Sorter100|8950_  = \new_Sorter100|8849_  | \new_Sorter100|8850_ ;
  assign \new_Sorter100|8951_  = \new_Sorter100|8851_  & \new_Sorter100|8852_ ;
  assign \new_Sorter100|8952_  = \new_Sorter100|8851_  | \new_Sorter100|8852_ ;
  assign \new_Sorter100|8953_  = \new_Sorter100|8853_  & \new_Sorter100|8854_ ;
  assign \new_Sorter100|8954_  = \new_Sorter100|8853_  | \new_Sorter100|8854_ ;
  assign \new_Sorter100|8955_  = \new_Sorter100|8855_  & \new_Sorter100|8856_ ;
  assign \new_Sorter100|8956_  = \new_Sorter100|8855_  | \new_Sorter100|8856_ ;
  assign \new_Sorter100|8957_  = \new_Sorter100|8857_  & \new_Sorter100|8858_ ;
  assign \new_Sorter100|8958_  = \new_Sorter100|8857_  | \new_Sorter100|8858_ ;
  assign \new_Sorter100|8959_  = \new_Sorter100|8859_  & \new_Sorter100|8860_ ;
  assign \new_Sorter100|8960_  = \new_Sorter100|8859_  | \new_Sorter100|8860_ ;
  assign \new_Sorter100|8961_  = \new_Sorter100|8861_  & \new_Sorter100|8862_ ;
  assign \new_Sorter100|8962_  = \new_Sorter100|8861_  | \new_Sorter100|8862_ ;
  assign \new_Sorter100|8963_  = \new_Sorter100|8863_  & \new_Sorter100|8864_ ;
  assign \new_Sorter100|8964_  = \new_Sorter100|8863_  | \new_Sorter100|8864_ ;
  assign \new_Sorter100|8965_  = \new_Sorter100|8865_  & \new_Sorter100|8866_ ;
  assign \new_Sorter100|8966_  = \new_Sorter100|8865_  | \new_Sorter100|8866_ ;
  assign \new_Sorter100|8967_  = \new_Sorter100|8867_  & \new_Sorter100|8868_ ;
  assign \new_Sorter100|8968_  = \new_Sorter100|8867_  | \new_Sorter100|8868_ ;
  assign \new_Sorter100|8969_  = \new_Sorter100|8869_  & \new_Sorter100|8870_ ;
  assign \new_Sorter100|8970_  = \new_Sorter100|8869_  | \new_Sorter100|8870_ ;
  assign \new_Sorter100|8971_  = \new_Sorter100|8871_  & \new_Sorter100|8872_ ;
  assign \new_Sorter100|8972_  = \new_Sorter100|8871_  | \new_Sorter100|8872_ ;
  assign \new_Sorter100|8973_  = \new_Sorter100|8873_  & \new_Sorter100|8874_ ;
  assign \new_Sorter100|8974_  = \new_Sorter100|8873_  | \new_Sorter100|8874_ ;
  assign \new_Sorter100|8975_  = \new_Sorter100|8875_  & \new_Sorter100|8876_ ;
  assign \new_Sorter100|8976_  = \new_Sorter100|8875_  | \new_Sorter100|8876_ ;
  assign \new_Sorter100|8977_  = \new_Sorter100|8877_  & \new_Sorter100|8878_ ;
  assign \new_Sorter100|8978_  = \new_Sorter100|8877_  | \new_Sorter100|8878_ ;
  assign \new_Sorter100|8979_  = \new_Sorter100|8879_  & \new_Sorter100|8880_ ;
  assign \new_Sorter100|8980_  = \new_Sorter100|8879_  | \new_Sorter100|8880_ ;
  assign \new_Sorter100|8981_  = \new_Sorter100|8881_  & \new_Sorter100|8882_ ;
  assign \new_Sorter100|8982_  = \new_Sorter100|8881_  | \new_Sorter100|8882_ ;
  assign \new_Sorter100|8983_  = \new_Sorter100|8883_  & \new_Sorter100|8884_ ;
  assign \new_Sorter100|8984_  = \new_Sorter100|8883_  | \new_Sorter100|8884_ ;
  assign \new_Sorter100|8985_  = \new_Sorter100|8885_  & \new_Sorter100|8886_ ;
  assign \new_Sorter100|8986_  = \new_Sorter100|8885_  | \new_Sorter100|8886_ ;
  assign \new_Sorter100|8987_  = \new_Sorter100|8887_  & \new_Sorter100|8888_ ;
  assign \new_Sorter100|8988_  = \new_Sorter100|8887_  | \new_Sorter100|8888_ ;
  assign \new_Sorter100|8989_  = \new_Sorter100|8889_  & \new_Sorter100|8890_ ;
  assign \new_Sorter100|8990_  = \new_Sorter100|8889_  | \new_Sorter100|8890_ ;
  assign \new_Sorter100|8991_  = \new_Sorter100|8891_  & \new_Sorter100|8892_ ;
  assign \new_Sorter100|8992_  = \new_Sorter100|8891_  | \new_Sorter100|8892_ ;
  assign \new_Sorter100|8993_  = \new_Sorter100|8893_  & \new_Sorter100|8894_ ;
  assign \new_Sorter100|8994_  = \new_Sorter100|8893_  | \new_Sorter100|8894_ ;
  assign \new_Sorter100|8995_  = \new_Sorter100|8895_  & \new_Sorter100|8896_ ;
  assign \new_Sorter100|8996_  = \new_Sorter100|8895_  | \new_Sorter100|8896_ ;
  assign \new_Sorter100|8997_  = \new_Sorter100|8897_  & \new_Sorter100|8898_ ;
  assign \new_Sorter100|8998_  = \new_Sorter100|8897_  | \new_Sorter100|8898_ ;
  assign \new_Sorter100|9000_  = \new_Sorter100|8900_  & \new_Sorter100|8901_ ;
  assign \new_Sorter100|9001_  = \new_Sorter100|8900_  | \new_Sorter100|8901_ ;
  assign \new_Sorter100|9002_  = \new_Sorter100|8902_  & \new_Sorter100|8903_ ;
  assign \new_Sorter100|9003_  = \new_Sorter100|8902_  | \new_Sorter100|8903_ ;
  assign \new_Sorter100|9004_  = \new_Sorter100|8904_  & \new_Sorter100|8905_ ;
  assign \new_Sorter100|9005_  = \new_Sorter100|8904_  | \new_Sorter100|8905_ ;
  assign \new_Sorter100|9006_  = \new_Sorter100|8906_  & \new_Sorter100|8907_ ;
  assign \new_Sorter100|9007_  = \new_Sorter100|8906_  | \new_Sorter100|8907_ ;
  assign \new_Sorter100|9008_  = \new_Sorter100|8908_  & \new_Sorter100|8909_ ;
  assign \new_Sorter100|9009_  = \new_Sorter100|8908_  | \new_Sorter100|8909_ ;
  assign \new_Sorter100|9010_  = \new_Sorter100|8910_  & \new_Sorter100|8911_ ;
  assign \new_Sorter100|9011_  = \new_Sorter100|8910_  | \new_Sorter100|8911_ ;
  assign \new_Sorter100|9012_  = \new_Sorter100|8912_  & \new_Sorter100|8913_ ;
  assign \new_Sorter100|9013_  = \new_Sorter100|8912_  | \new_Sorter100|8913_ ;
  assign \new_Sorter100|9014_  = \new_Sorter100|8914_  & \new_Sorter100|8915_ ;
  assign \new_Sorter100|9015_  = \new_Sorter100|8914_  | \new_Sorter100|8915_ ;
  assign \new_Sorter100|9016_  = \new_Sorter100|8916_  & \new_Sorter100|8917_ ;
  assign \new_Sorter100|9017_  = \new_Sorter100|8916_  | \new_Sorter100|8917_ ;
  assign \new_Sorter100|9018_  = \new_Sorter100|8918_  & \new_Sorter100|8919_ ;
  assign \new_Sorter100|9019_  = \new_Sorter100|8918_  | \new_Sorter100|8919_ ;
  assign \new_Sorter100|9020_  = \new_Sorter100|8920_  & \new_Sorter100|8921_ ;
  assign \new_Sorter100|9021_  = \new_Sorter100|8920_  | \new_Sorter100|8921_ ;
  assign \new_Sorter100|9022_  = \new_Sorter100|8922_  & \new_Sorter100|8923_ ;
  assign \new_Sorter100|9023_  = \new_Sorter100|8922_  | \new_Sorter100|8923_ ;
  assign \new_Sorter100|9024_  = \new_Sorter100|8924_  & \new_Sorter100|8925_ ;
  assign \new_Sorter100|9025_  = \new_Sorter100|8924_  | \new_Sorter100|8925_ ;
  assign \new_Sorter100|9026_  = \new_Sorter100|8926_  & \new_Sorter100|8927_ ;
  assign \new_Sorter100|9027_  = \new_Sorter100|8926_  | \new_Sorter100|8927_ ;
  assign \new_Sorter100|9028_  = \new_Sorter100|8928_  & \new_Sorter100|8929_ ;
  assign \new_Sorter100|9029_  = \new_Sorter100|8928_  | \new_Sorter100|8929_ ;
  assign \new_Sorter100|9030_  = \new_Sorter100|8930_  & \new_Sorter100|8931_ ;
  assign \new_Sorter100|9031_  = \new_Sorter100|8930_  | \new_Sorter100|8931_ ;
  assign \new_Sorter100|9032_  = \new_Sorter100|8932_  & \new_Sorter100|8933_ ;
  assign \new_Sorter100|9033_  = \new_Sorter100|8932_  | \new_Sorter100|8933_ ;
  assign \new_Sorter100|9034_  = \new_Sorter100|8934_  & \new_Sorter100|8935_ ;
  assign \new_Sorter100|9035_  = \new_Sorter100|8934_  | \new_Sorter100|8935_ ;
  assign \new_Sorter100|9036_  = \new_Sorter100|8936_  & \new_Sorter100|8937_ ;
  assign \new_Sorter100|9037_  = \new_Sorter100|8936_  | \new_Sorter100|8937_ ;
  assign \new_Sorter100|9038_  = \new_Sorter100|8938_  & \new_Sorter100|8939_ ;
  assign \new_Sorter100|9039_  = \new_Sorter100|8938_  | \new_Sorter100|8939_ ;
  assign \new_Sorter100|9040_  = \new_Sorter100|8940_  & \new_Sorter100|8941_ ;
  assign \new_Sorter100|9041_  = \new_Sorter100|8940_  | \new_Sorter100|8941_ ;
  assign \new_Sorter100|9042_  = \new_Sorter100|8942_  & \new_Sorter100|8943_ ;
  assign \new_Sorter100|9043_  = \new_Sorter100|8942_  | \new_Sorter100|8943_ ;
  assign \new_Sorter100|9044_  = \new_Sorter100|8944_  & \new_Sorter100|8945_ ;
  assign \new_Sorter100|9045_  = \new_Sorter100|8944_  | \new_Sorter100|8945_ ;
  assign \new_Sorter100|9046_  = \new_Sorter100|8946_  & \new_Sorter100|8947_ ;
  assign \new_Sorter100|9047_  = \new_Sorter100|8946_  | \new_Sorter100|8947_ ;
  assign \new_Sorter100|9048_  = \new_Sorter100|8948_  & \new_Sorter100|8949_ ;
  assign \new_Sorter100|9049_  = \new_Sorter100|8948_  | \new_Sorter100|8949_ ;
  assign \new_Sorter100|9050_  = \new_Sorter100|8950_  & \new_Sorter100|8951_ ;
  assign \new_Sorter100|9051_  = \new_Sorter100|8950_  | \new_Sorter100|8951_ ;
  assign \new_Sorter100|9052_  = \new_Sorter100|8952_  & \new_Sorter100|8953_ ;
  assign \new_Sorter100|9053_  = \new_Sorter100|8952_  | \new_Sorter100|8953_ ;
  assign \new_Sorter100|9054_  = \new_Sorter100|8954_  & \new_Sorter100|8955_ ;
  assign \new_Sorter100|9055_  = \new_Sorter100|8954_  | \new_Sorter100|8955_ ;
  assign \new_Sorter100|9056_  = \new_Sorter100|8956_  & \new_Sorter100|8957_ ;
  assign \new_Sorter100|9057_  = \new_Sorter100|8956_  | \new_Sorter100|8957_ ;
  assign \new_Sorter100|9058_  = \new_Sorter100|8958_  & \new_Sorter100|8959_ ;
  assign \new_Sorter100|9059_  = \new_Sorter100|8958_  | \new_Sorter100|8959_ ;
  assign \new_Sorter100|9060_  = \new_Sorter100|8960_  & \new_Sorter100|8961_ ;
  assign \new_Sorter100|9061_  = \new_Sorter100|8960_  | \new_Sorter100|8961_ ;
  assign \new_Sorter100|9062_  = \new_Sorter100|8962_  & \new_Sorter100|8963_ ;
  assign \new_Sorter100|9063_  = \new_Sorter100|8962_  | \new_Sorter100|8963_ ;
  assign \new_Sorter100|9064_  = \new_Sorter100|8964_  & \new_Sorter100|8965_ ;
  assign \new_Sorter100|9065_  = \new_Sorter100|8964_  | \new_Sorter100|8965_ ;
  assign \new_Sorter100|9066_  = \new_Sorter100|8966_  & \new_Sorter100|8967_ ;
  assign \new_Sorter100|9067_  = \new_Sorter100|8966_  | \new_Sorter100|8967_ ;
  assign \new_Sorter100|9068_  = \new_Sorter100|8968_  & \new_Sorter100|8969_ ;
  assign \new_Sorter100|9069_  = \new_Sorter100|8968_  | \new_Sorter100|8969_ ;
  assign \new_Sorter100|9070_  = \new_Sorter100|8970_  & \new_Sorter100|8971_ ;
  assign \new_Sorter100|9071_  = \new_Sorter100|8970_  | \new_Sorter100|8971_ ;
  assign \new_Sorter100|9072_  = \new_Sorter100|8972_  & \new_Sorter100|8973_ ;
  assign \new_Sorter100|9073_  = \new_Sorter100|8972_  | \new_Sorter100|8973_ ;
  assign \new_Sorter100|9074_  = \new_Sorter100|8974_  & \new_Sorter100|8975_ ;
  assign \new_Sorter100|9075_  = \new_Sorter100|8974_  | \new_Sorter100|8975_ ;
  assign \new_Sorter100|9076_  = \new_Sorter100|8976_  & \new_Sorter100|8977_ ;
  assign \new_Sorter100|9077_  = \new_Sorter100|8976_  | \new_Sorter100|8977_ ;
  assign \new_Sorter100|9078_  = \new_Sorter100|8978_  & \new_Sorter100|8979_ ;
  assign \new_Sorter100|9079_  = \new_Sorter100|8978_  | \new_Sorter100|8979_ ;
  assign \new_Sorter100|9080_  = \new_Sorter100|8980_  & \new_Sorter100|8981_ ;
  assign \new_Sorter100|9081_  = \new_Sorter100|8980_  | \new_Sorter100|8981_ ;
  assign \new_Sorter100|9082_  = \new_Sorter100|8982_  & \new_Sorter100|8983_ ;
  assign \new_Sorter100|9083_  = \new_Sorter100|8982_  | \new_Sorter100|8983_ ;
  assign \new_Sorter100|9084_  = \new_Sorter100|8984_  & \new_Sorter100|8985_ ;
  assign \new_Sorter100|9085_  = \new_Sorter100|8984_  | \new_Sorter100|8985_ ;
  assign \new_Sorter100|9086_  = \new_Sorter100|8986_  & \new_Sorter100|8987_ ;
  assign \new_Sorter100|9087_  = \new_Sorter100|8986_  | \new_Sorter100|8987_ ;
  assign \new_Sorter100|9088_  = \new_Sorter100|8988_  & \new_Sorter100|8989_ ;
  assign \new_Sorter100|9089_  = \new_Sorter100|8988_  | \new_Sorter100|8989_ ;
  assign \new_Sorter100|9090_  = \new_Sorter100|8990_  & \new_Sorter100|8991_ ;
  assign \new_Sorter100|9091_  = \new_Sorter100|8990_  | \new_Sorter100|8991_ ;
  assign \new_Sorter100|9092_  = \new_Sorter100|8992_  & \new_Sorter100|8993_ ;
  assign \new_Sorter100|9093_  = \new_Sorter100|8992_  | \new_Sorter100|8993_ ;
  assign \new_Sorter100|9094_  = \new_Sorter100|8994_  & \new_Sorter100|8995_ ;
  assign \new_Sorter100|9095_  = \new_Sorter100|8994_  | \new_Sorter100|8995_ ;
  assign \new_Sorter100|9096_  = \new_Sorter100|8996_  & \new_Sorter100|8997_ ;
  assign \new_Sorter100|9097_  = \new_Sorter100|8996_  | \new_Sorter100|8997_ ;
  assign \new_Sorter100|9098_  = \new_Sorter100|8998_  & \new_Sorter100|8999_ ;
  assign \new_Sorter100|9099_  = \new_Sorter100|8998_  | \new_Sorter100|8999_ ;
  assign \new_Sorter100|9100_  = \new_Sorter100|9000_ ;
  assign \new_Sorter100|9199_  = \new_Sorter100|9099_ ;
  assign \new_Sorter100|9101_  = \new_Sorter100|9001_  & \new_Sorter100|9002_ ;
  assign \new_Sorter100|9102_  = \new_Sorter100|9001_  | \new_Sorter100|9002_ ;
  assign \new_Sorter100|9103_  = \new_Sorter100|9003_  & \new_Sorter100|9004_ ;
  assign \new_Sorter100|9104_  = \new_Sorter100|9003_  | \new_Sorter100|9004_ ;
  assign \new_Sorter100|9105_  = \new_Sorter100|9005_  & \new_Sorter100|9006_ ;
  assign \new_Sorter100|9106_  = \new_Sorter100|9005_  | \new_Sorter100|9006_ ;
  assign \new_Sorter100|9107_  = \new_Sorter100|9007_  & \new_Sorter100|9008_ ;
  assign \new_Sorter100|9108_  = \new_Sorter100|9007_  | \new_Sorter100|9008_ ;
  assign \new_Sorter100|9109_  = \new_Sorter100|9009_  & \new_Sorter100|9010_ ;
  assign \new_Sorter100|9110_  = \new_Sorter100|9009_  | \new_Sorter100|9010_ ;
  assign \new_Sorter100|9111_  = \new_Sorter100|9011_  & \new_Sorter100|9012_ ;
  assign \new_Sorter100|9112_  = \new_Sorter100|9011_  | \new_Sorter100|9012_ ;
  assign \new_Sorter100|9113_  = \new_Sorter100|9013_  & \new_Sorter100|9014_ ;
  assign \new_Sorter100|9114_  = \new_Sorter100|9013_  | \new_Sorter100|9014_ ;
  assign \new_Sorter100|9115_  = \new_Sorter100|9015_  & \new_Sorter100|9016_ ;
  assign \new_Sorter100|9116_  = \new_Sorter100|9015_  | \new_Sorter100|9016_ ;
  assign \new_Sorter100|9117_  = \new_Sorter100|9017_  & \new_Sorter100|9018_ ;
  assign \new_Sorter100|9118_  = \new_Sorter100|9017_  | \new_Sorter100|9018_ ;
  assign \new_Sorter100|9119_  = \new_Sorter100|9019_  & \new_Sorter100|9020_ ;
  assign \new_Sorter100|9120_  = \new_Sorter100|9019_  | \new_Sorter100|9020_ ;
  assign \new_Sorter100|9121_  = \new_Sorter100|9021_  & \new_Sorter100|9022_ ;
  assign \new_Sorter100|9122_  = \new_Sorter100|9021_  | \new_Sorter100|9022_ ;
  assign \new_Sorter100|9123_  = \new_Sorter100|9023_  & \new_Sorter100|9024_ ;
  assign \new_Sorter100|9124_  = \new_Sorter100|9023_  | \new_Sorter100|9024_ ;
  assign \new_Sorter100|9125_  = \new_Sorter100|9025_  & \new_Sorter100|9026_ ;
  assign \new_Sorter100|9126_  = \new_Sorter100|9025_  | \new_Sorter100|9026_ ;
  assign \new_Sorter100|9127_  = \new_Sorter100|9027_  & \new_Sorter100|9028_ ;
  assign \new_Sorter100|9128_  = \new_Sorter100|9027_  | \new_Sorter100|9028_ ;
  assign \new_Sorter100|9129_  = \new_Sorter100|9029_  & \new_Sorter100|9030_ ;
  assign \new_Sorter100|9130_  = \new_Sorter100|9029_  | \new_Sorter100|9030_ ;
  assign \new_Sorter100|9131_  = \new_Sorter100|9031_  & \new_Sorter100|9032_ ;
  assign \new_Sorter100|9132_  = \new_Sorter100|9031_  | \new_Sorter100|9032_ ;
  assign \new_Sorter100|9133_  = \new_Sorter100|9033_  & \new_Sorter100|9034_ ;
  assign \new_Sorter100|9134_  = \new_Sorter100|9033_  | \new_Sorter100|9034_ ;
  assign \new_Sorter100|9135_  = \new_Sorter100|9035_  & \new_Sorter100|9036_ ;
  assign \new_Sorter100|9136_  = \new_Sorter100|9035_  | \new_Sorter100|9036_ ;
  assign \new_Sorter100|9137_  = \new_Sorter100|9037_  & \new_Sorter100|9038_ ;
  assign \new_Sorter100|9138_  = \new_Sorter100|9037_  | \new_Sorter100|9038_ ;
  assign \new_Sorter100|9139_  = \new_Sorter100|9039_  & \new_Sorter100|9040_ ;
  assign \new_Sorter100|9140_  = \new_Sorter100|9039_  | \new_Sorter100|9040_ ;
  assign \new_Sorter100|9141_  = \new_Sorter100|9041_  & \new_Sorter100|9042_ ;
  assign \new_Sorter100|9142_  = \new_Sorter100|9041_  | \new_Sorter100|9042_ ;
  assign \new_Sorter100|9143_  = \new_Sorter100|9043_  & \new_Sorter100|9044_ ;
  assign \new_Sorter100|9144_  = \new_Sorter100|9043_  | \new_Sorter100|9044_ ;
  assign \new_Sorter100|9145_  = \new_Sorter100|9045_  & \new_Sorter100|9046_ ;
  assign \new_Sorter100|9146_  = \new_Sorter100|9045_  | \new_Sorter100|9046_ ;
  assign \new_Sorter100|9147_  = \new_Sorter100|9047_  & \new_Sorter100|9048_ ;
  assign \new_Sorter100|9148_  = \new_Sorter100|9047_  | \new_Sorter100|9048_ ;
  assign \new_Sorter100|9149_  = \new_Sorter100|9049_  & \new_Sorter100|9050_ ;
  assign \new_Sorter100|9150_  = \new_Sorter100|9049_  | \new_Sorter100|9050_ ;
  assign \new_Sorter100|9151_  = \new_Sorter100|9051_  & \new_Sorter100|9052_ ;
  assign \new_Sorter100|9152_  = \new_Sorter100|9051_  | \new_Sorter100|9052_ ;
  assign \new_Sorter100|9153_  = \new_Sorter100|9053_  & \new_Sorter100|9054_ ;
  assign \new_Sorter100|9154_  = \new_Sorter100|9053_  | \new_Sorter100|9054_ ;
  assign \new_Sorter100|9155_  = \new_Sorter100|9055_  & \new_Sorter100|9056_ ;
  assign \new_Sorter100|9156_  = \new_Sorter100|9055_  | \new_Sorter100|9056_ ;
  assign \new_Sorter100|9157_  = \new_Sorter100|9057_  & \new_Sorter100|9058_ ;
  assign \new_Sorter100|9158_  = \new_Sorter100|9057_  | \new_Sorter100|9058_ ;
  assign \new_Sorter100|9159_  = \new_Sorter100|9059_  & \new_Sorter100|9060_ ;
  assign \new_Sorter100|9160_  = \new_Sorter100|9059_  | \new_Sorter100|9060_ ;
  assign \new_Sorter100|9161_  = \new_Sorter100|9061_  & \new_Sorter100|9062_ ;
  assign \new_Sorter100|9162_  = \new_Sorter100|9061_  | \new_Sorter100|9062_ ;
  assign \new_Sorter100|9163_  = \new_Sorter100|9063_  & \new_Sorter100|9064_ ;
  assign \new_Sorter100|9164_  = \new_Sorter100|9063_  | \new_Sorter100|9064_ ;
  assign \new_Sorter100|9165_  = \new_Sorter100|9065_  & \new_Sorter100|9066_ ;
  assign \new_Sorter100|9166_  = \new_Sorter100|9065_  | \new_Sorter100|9066_ ;
  assign \new_Sorter100|9167_  = \new_Sorter100|9067_  & \new_Sorter100|9068_ ;
  assign \new_Sorter100|9168_  = \new_Sorter100|9067_  | \new_Sorter100|9068_ ;
  assign \new_Sorter100|9169_  = \new_Sorter100|9069_  & \new_Sorter100|9070_ ;
  assign \new_Sorter100|9170_  = \new_Sorter100|9069_  | \new_Sorter100|9070_ ;
  assign \new_Sorter100|9171_  = \new_Sorter100|9071_  & \new_Sorter100|9072_ ;
  assign \new_Sorter100|9172_  = \new_Sorter100|9071_  | \new_Sorter100|9072_ ;
  assign \new_Sorter100|9173_  = \new_Sorter100|9073_  & \new_Sorter100|9074_ ;
  assign \new_Sorter100|9174_  = \new_Sorter100|9073_  | \new_Sorter100|9074_ ;
  assign \new_Sorter100|9175_  = \new_Sorter100|9075_  & \new_Sorter100|9076_ ;
  assign \new_Sorter100|9176_  = \new_Sorter100|9075_  | \new_Sorter100|9076_ ;
  assign \new_Sorter100|9177_  = \new_Sorter100|9077_  & \new_Sorter100|9078_ ;
  assign \new_Sorter100|9178_  = \new_Sorter100|9077_  | \new_Sorter100|9078_ ;
  assign \new_Sorter100|9179_  = \new_Sorter100|9079_  & \new_Sorter100|9080_ ;
  assign \new_Sorter100|9180_  = \new_Sorter100|9079_  | \new_Sorter100|9080_ ;
  assign \new_Sorter100|9181_  = \new_Sorter100|9081_  & \new_Sorter100|9082_ ;
  assign \new_Sorter100|9182_  = \new_Sorter100|9081_  | \new_Sorter100|9082_ ;
  assign \new_Sorter100|9183_  = \new_Sorter100|9083_  & \new_Sorter100|9084_ ;
  assign \new_Sorter100|9184_  = \new_Sorter100|9083_  | \new_Sorter100|9084_ ;
  assign \new_Sorter100|9185_  = \new_Sorter100|9085_  & \new_Sorter100|9086_ ;
  assign \new_Sorter100|9186_  = \new_Sorter100|9085_  | \new_Sorter100|9086_ ;
  assign \new_Sorter100|9187_  = \new_Sorter100|9087_  & \new_Sorter100|9088_ ;
  assign \new_Sorter100|9188_  = \new_Sorter100|9087_  | \new_Sorter100|9088_ ;
  assign \new_Sorter100|9189_  = \new_Sorter100|9089_  & \new_Sorter100|9090_ ;
  assign \new_Sorter100|9190_  = \new_Sorter100|9089_  | \new_Sorter100|9090_ ;
  assign \new_Sorter100|9191_  = \new_Sorter100|9091_  & \new_Sorter100|9092_ ;
  assign \new_Sorter100|9192_  = \new_Sorter100|9091_  | \new_Sorter100|9092_ ;
  assign \new_Sorter100|9193_  = \new_Sorter100|9093_  & \new_Sorter100|9094_ ;
  assign \new_Sorter100|9194_  = \new_Sorter100|9093_  | \new_Sorter100|9094_ ;
  assign \new_Sorter100|9195_  = \new_Sorter100|9095_  & \new_Sorter100|9096_ ;
  assign \new_Sorter100|9196_  = \new_Sorter100|9095_  | \new_Sorter100|9096_ ;
  assign \new_Sorter100|9197_  = \new_Sorter100|9097_  & \new_Sorter100|9098_ ;
  assign \new_Sorter100|9198_  = \new_Sorter100|9097_  | \new_Sorter100|9098_ ;
  assign \new_Sorter100|9200_  = \new_Sorter100|9100_  & \new_Sorter100|9101_ ;
  assign \new_Sorter100|9201_  = \new_Sorter100|9100_  | \new_Sorter100|9101_ ;
  assign \new_Sorter100|9202_  = \new_Sorter100|9102_  & \new_Sorter100|9103_ ;
  assign \new_Sorter100|9203_  = \new_Sorter100|9102_  | \new_Sorter100|9103_ ;
  assign \new_Sorter100|9204_  = \new_Sorter100|9104_  & \new_Sorter100|9105_ ;
  assign \new_Sorter100|9205_  = \new_Sorter100|9104_  | \new_Sorter100|9105_ ;
  assign \new_Sorter100|9206_  = \new_Sorter100|9106_  & \new_Sorter100|9107_ ;
  assign \new_Sorter100|9207_  = \new_Sorter100|9106_  | \new_Sorter100|9107_ ;
  assign \new_Sorter100|9208_  = \new_Sorter100|9108_  & \new_Sorter100|9109_ ;
  assign \new_Sorter100|9209_  = \new_Sorter100|9108_  | \new_Sorter100|9109_ ;
  assign \new_Sorter100|9210_  = \new_Sorter100|9110_  & \new_Sorter100|9111_ ;
  assign \new_Sorter100|9211_  = \new_Sorter100|9110_  | \new_Sorter100|9111_ ;
  assign \new_Sorter100|9212_  = \new_Sorter100|9112_  & \new_Sorter100|9113_ ;
  assign \new_Sorter100|9213_  = \new_Sorter100|9112_  | \new_Sorter100|9113_ ;
  assign \new_Sorter100|9214_  = \new_Sorter100|9114_  & \new_Sorter100|9115_ ;
  assign \new_Sorter100|9215_  = \new_Sorter100|9114_  | \new_Sorter100|9115_ ;
  assign \new_Sorter100|9216_  = \new_Sorter100|9116_  & \new_Sorter100|9117_ ;
  assign \new_Sorter100|9217_  = \new_Sorter100|9116_  | \new_Sorter100|9117_ ;
  assign \new_Sorter100|9218_  = \new_Sorter100|9118_  & \new_Sorter100|9119_ ;
  assign \new_Sorter100|9219_  = \new_Sorter100|9118_  | \new_Sorter100|9119_ ;
  assign \new_Sorter100|9220_  = \new_Sorter100|9120_  & \new_Sorter100|9121_ ;
  assign \new_Sorter100|9221_  = \new_Sorter100|9120_  | \new_Sorter100|9121_ ;
  assign \new_Sorter100|9222_  = \new_Sorter100|9122_  & \new_Sorter100|9123_ ;
  assign \new_Sorter100|9223_  = \new_Sorter100|9122_  | \new_Sorter100|9123_ ;
  assign \new_Sorter100|9224_  = \new_Sorter100|9124_  & \new_Sorter100|9125_ ;
  assign \new_Sorter100|9225_  = \new_Sorter100|9124_  | \new_Sorter100|9125_ ;
  assign \new_Sorter100|9226_  = \new_Sorter100|9126_  & \new_Sorter100|9127_ ;
  assign \new_Sorter100|9227_  = \new_Sorter100|9126_  | \new_Sorter100|9127_ ;
  assign \new_Sorter100|9228_  = \new_Sorter100|9128_  & \new_Sorter100|9129_ ;
  assign \new_Sorter100|9229_  = \new_Sorter100|9128_  | \new_Sorter100|9129_ ;
  assign \new_Sorter100|9230_  = \new_Sorter100|9130_  & \new_Sorter100|9131_ ;
  assign \new_Sorter100|9231_  = \new_Sorter100|9130_  | \new_Sorter100|9131_ ;
  assign \new_Sorter100|9232_  = \new_Sorter100|9132_  & \new_Sorter100|9133_ ;
  assign \new_Sorter100|9233_  = \new_Sorter100|9132_  | \new_Sorter100|9133_ ;
  assign \new_Sorter100|9234_  = \new_Sorter100|9134_  & \new_Sorter100|9135_ ;
  assign \new_Sorter100|9235_  = \new_Sorter100|9134_  | \new_Sorter100|9135_ ;
  assign \new_Sorter100|9236_  = \new_Sorter100|9136_  & \new_Sorter100|9137_ ;
  assign \new_Sorter100|9237_  = \new_Sorter100|9136_  | \new_Sorter100|9137_ ;
  assign \new_Sorter100|9238_  = \new_Sorter100|9138_  & \new_Sorter100|9139_ ;
  assign \new_Sorter100|9239_  = \new_Sorter100|9138_  | \new_Sorter100|9139_ ;
  assign \new_Sorter100|9240_  = \new_Sorter100|9140_  & \new_Sorter100|9141_ ;
  assign \new_Sorter100|9241_  = \new_Sorter100|9140_  | \new_Sorter100|9141_ ;
  assign \new_Sorter100|9242_  = \new_Sorter100|9142_  & \new_Sorter100|9143_ ;
  assign \new_Sorter100|9243_  = \new_Sorter100|9142_  | \new_Sorter100|9143_ ;
  assign \new_Sorter100|9244_  = \new_Sorter100|9144_  & \new_Sorter100|9145_ ;
  assign \new_Sorter100|9245_  = \new_Sorter100|9144_  | \new_Sorter100|9145_ ;
  assign \new_Sorter100|9246_  = \new_Sorter100|9146_  & \new_Sorter100|9147_ ;
  assign \new_Sorter100|9247_  = \new_Sorter100|9146_  | \new_Sorter100|9147_ ;
  assign \new_Sorter100|9248_  = \new_Sorter100|9148_  & \new_Sorter100|9149_ ;
  assign \new_Sorter100|9249_  = \new_Sorter100|9148_  | \new_Sorter100|9149_ ;
  assign \new_Sorter100|9250_  = \new_Sorter100|9150_  & \new_Sorter100|9151_ ;
  assign \new_Sorter100|9251_  = \new_Sorter100|9150_  | \new_Sorter100|9151_ ;
  assign \new_Sorter100|9252_  = \new_Sorter100|9152_  & \new_Sorter100|9153_ ;
  assign \new_Sorter100|9253_  = \new_Sorter100|9152_  | \new_Sorter100|9153_ ;
  assign \new_Sorter100|9254_  = \new_Sorter100|9154_  & \new_Sorter100|9155_ ;
  assign \new_Sorter100|9255_  = \new_Sorter100|9154_  | \new_Sorter100|9155_ ;
  assign \new_Sorter100|9256_  = \new_Sorter100|9156_  & \new_Sorter100|9157_ ;
  assign \new_Sorter100|9257_  = \new_Sorter100|9156_  | \new_Sorter100|9157_ ;
  assign \new_Sorter100|9258_  = \new_Sorter100|9158_  & \new_Sorter100|9159_ ;
  assign \new_Sorter100|9259_  = \new_Sorter100|9158_  | \new_Sorter100|9159_ ;
  assign \new_Sorter100|9260_  = \new_Sorter100|9160_  & \new_Sorter100|9161_ ;
  assign \new_Sorter100|9261_  = \new_Sorter100|9160_  | \new_Sorter100|9161_ ;
  assign \new_Sorter100|9262_  = \new_Sorter100|9162_  & \new_Sorter100|9163_ ;
  assign \new_Sorter100|9263_  = \new_Sorter100|9162_  | \new_Sorter100|9163_ ;
  assign \new_Sorter100|9264_  = \new_Sorter100|9164_  & \new_Sorter100|9165_ ;
  assign \new_Sorter100|9265_  = \new_Sorter100|9164_  | \new_Sorter100|9165_ ;
  assign \new_Sorter100|9266_  = \new_Sorter100|9166_  & \new_Sorter100|9167_ ;
  assign \new_Sorter100|9267_  = \new_Sorter100|9166_  | \new_Sorter100|9167_ ;
  assign \new_Sorter100|9268_  = \new_Sorter100|9168_  & \new_Sorter100|9169_ ;
  assign \new_Sorter100|9269_  = \new_Sorter100|9168_  | \new_Sorter100|9169_ ;
  assign \new_Sorter100|9270_  = \new_Sorter100|9170_  & \new_Sorter100|9171_ ;
  assign \new_Sorter100|9271_  = \new_Sorter100|9170_  | \new_Sorter100|9171_ ;
  assign \new_Sorter100|9272_  = \new_Sorter100|9172_  & \new_Sorter100|9173_ ;
  assign \new_Sorter100|9273_  = \new_Sorter100|9172_  | \new_Sorter100|9173_ ;
  assign \new_Sorter100|9274_  = \new_Sorter100|9174_  & \new_Sorter100|9175_ ;
  assign \new_Sorter100|9275_  = \new_Sorter100|9174_  | \new_Sorter100|9175_ ;
  assign \new_Sorter100|9276_  = \new_Sorter100|9176_  & \new_Sorter100|9177_ ;
  assign \new_Sorter100|9277_  = \new_Sorter100|9176_  | \new_Sorter100|9177_ ;
  assign \new_Sorter100|9278_  = \new_Sorter100|9178_  & \new_Sorter100|9179_ ;
  assign \new_Sorter100|9279_  = \new_Sorter100|9178_  | \new_Sorter100|9179_ ;
  assign \new_Sorter100|9280_  = \new_Sorter100|9180_  & \new_Sorter100|9181_ ;
  assign \new_Sorter100|9281_  = \new_Sorter100|9180_  | \new_Sorter100|9181_ ;
  assign \new_Sorter100|9282_  = \new_Sorter100|9182_  & \new_Sorter100|9183_ ;
  assign \new_Sorter100|9283_  = \new_Sorter100|9182_  | \new_Sorter100|9183_ ;
  assign \new_Sorter100|9284_  = \new_Sorter100|9184_  & \new_Sorter100|9185_ ;
  assign \new_Sorter100|9285_  = \new_Sorter100|9184_  | \new_Sorter100|9185_ ;
  assign \new_Sorter100|9286_  = \new_Sorter100|9186_  & \new_Sorter100|9187_ ;
  assign \new_Sorter100|9287_  = \new_Sorter100|9186_  | \new_Sorter100|9187_ ;
  assign \new_Sorter100|9288_  = \new_Sorter100|9188_  & \new_Sorter100|9189_ ;
  assign \new_Sorter100|9289_  = \new_Sorter100|9188_  | \new_Sorter100|9189_ ;
  assign \new_Sorter100|9290_  = \new_Sorter100|9190_  & \new_Sorter100|9191_ ;
  assign \new_Sorter100|9291_  = \new_Sorter100|9190_  | \new_Sorter100|9191_ ;
  assign \new_Sorter100|9292_  = \new_Sorter100|9192_  & \new_Sorter100|9193_ ;
  assign \new_Sorter100|9293_  = \new_Sorter100|9192_  | \new_Sorter100|9193_ ;
  assign \new_Sorter100|9294_  = \new_Sorter100|9194_  & \new_Sorter100|9195_ ;
  assign \new_Sorter100|9295_  = \new_Sorter100|9194_  | \new_Sorter100|9195_ ;
  assign \new_Sorter100|9296_  = \new_Sorter100|9196_  & \new_Sorter100|9197_ ;
  assign \new_Sorter100|9297_  = \new_Sorter100|9196_  | \new_Sorter100|9197_ ;
  assign \new_Sorter100|9298_  = \new_Sorter100|9198_  & \new_Sorter100|9199_ ;
  assign \new_Sorter100|9299_  = \new_Sorter100|9198_  | \new_Sorter100|9199_ ;
  assign \new_Sorter100|9300_  = \new_Sorter100|9200_ ;
  assign \new_Sorter100|9399_  = \new_Sorter100|9299_ ;
  assign \new_Sorter100|9301_  = \new_Sorter100|9201_  & \new_Sorter100|9202_ ;
  assign \new_Sorter100|9302_  = \new_Sorter100|9201_  | \new_Sorter100|9202_ ;
  assign \new_Sorter100|9303_  = \new_Sorter100|9203_  & \new_Sorter100|9204_ ;
  assign \new_Sorter100|9304_  = \new_Sorter100|9203_  | \new_Sorter100|9204_ ;
  assign \new_Sorter100|9305_  = \new_Sorter100|9205_  & \new_Sorter100|9206_ ;
  assign \new_Sorter100|9306_  = \new_Sorter100|9205_  | \new_Sorter100|9206_ ;
  assign \new_Sorter100|9307_  = \new_Sorter100|9207_  & \new_Sorter100|9208_ ;
  assign \new_Sorter100|9308_  = \new_Sorter100|9207_  | \new_Sorter100|9208_ ;
  assign \new_Sorter100|9309_  = \new_Sorter100|9209_  & \new_Sorter100|9210_ ;
  assign \new_Sorter100|9310_  = \new_Sorter100|9209_  | \new_Sorter100|9210_ ;
  assign \new_Sorter100|9311_  = \new_Sorter100|9211_  & \new_Sorter100|9212_ ;
  assign \new_Sorter100|9312_  = \new_Sorter100|9211_  | \new_Sorter100|9212_ ;
  assign \new_Sorter100|9313_  = \new_Sorter100|9213_  & \new_Sorter100|9214_ ;
  assign \new_Sorter100|9314_  = \new_Sorter100|9213_  | \new_Sorter100|9214_ ;
  assign \new_Sorter100|9315_  = \new_Sorter100|9215_  & \new_Sorter100|9216_ ;
  assign \new_Sorter100|9316_  = \new_Sorter100|9215_  | \new_Sorter100|9216_ ;
  assign \new_Sorter100|9317_  = \new_Sorter100|9217_  & \new_Sorter100|9218_ ;
  assign \new_Sorter100|9318_  = \new_Sorter100|9217_  | \new_Sorter100|9218_ ;
  assign \new_Sorter100|9319_  = \new_Sorter100|9219_  & \new_Sorter100|9220_ ;
  assign \new_Sorter100|9320_  = \new_Sorter100|9219_  | \new_Sorter100|9220_ ;
  assign \new_Sorter100|9321_  = \new_Sorter100|9221_  & \new_Sorter100|9222_ ;
  assign \new_Sorter100|9322_  = \new_Sorter100|9221_  | \new_Sorter100|9222_ ;
  assign \new_Sorter100|9323_  = \new_Sorter100|9223_  & \new_Sorter100|9224_ ;
  assign \new_Sorter100|9324_  = \new_Sorter100|9223_  | \new_Sorter100|9224_ ;
  assign \new_Sorter100|9325_  = \new_Sorter100|9225_  & \new_Sorter100|9226_ ;
  assign \new_Sorter100|9326_  = \new_Sorter100|9225_  | \new_Sorter100|9226_ ;
  assign \new_Sorter100|9327_  = \new_Sorter100|9227_  & \new_Sorter100|9228_ ;
  assign \new_Sorter100|9328_  = \new_Sorter100|9227_  | \new_Sorter100|9228_ ;
  assign \new_Sorter100|9329_  = \new_Sorter100|9229_  & \new_Sorter100|9230_ ;
  assign \new_Sorter100|9330_  = \new_Sorter100|9229_  | \new_Sorter100|9230_ ;
  assign \new_Sorter100|9331_  = \new_Sorter100|9231_  & \new_Sorter100|9232_ ;
  assign \new_Sorter100|9332_  = \new_Sorter100|9231_  | \new_Sorter100|9232_ ;
  assign \new_Sorter100|9333_  = \new_Sorter100|9233_  & \new_Sorter100|9234_ ;
  assign \new_Sorter100|9334_  = \new_Sorter100|9233_  | \new_Sorter100|9234_ ;
  assign \new_Sorter100|9335_  = \new_Sorter100|9235_  & \new_Sorter100|9236_ ;
  assign \new_Sorter100|9336_  = \new_Sorter100|9235_  | \new_Sorter100|9236_ ;
  assign \new_Sorter100|9337_  = \new_Sorter100|9237_  & \new_Sorter100|9238_ ;
  assign \new_Sorter100|9338_  = \new_Sorter100|9237_  | \new_Sorter100|9238_ ;
  assign \new_Sorter100|9339_  = \new_Sorter100|9239_  & \new_Sorter100|9240_ ;
  assign \new_Sorter100|9340_  = \new_Sorter100|9239_  | \new_Sorter100|9240_ ;
  assign \new_Sorter100|9341_  = \new_Sorter100|9241_  & \new_Sorter100|9242_ ;
  assign \new_Sorter100|9342_  = \new_Sorter100|9241_  | \new_Sorter100|9242_ ;
  assign \new_Sorter100|9343_  = \new_Sorter100|9243_  & \new_Sorter100|9244_ ;
  assign \new_Sorter100|9344_  = \new_Sorter100|9243_  | \new_Sorter100|9244_ ;
  assign \new_Sorter100|9345_  = \new_Sorter100|9245_  & \new_Sorter100|9246_ ;
  assign \new_Sorter100|9346_  = \new_Sorter100|9245_  | \new_Sorter100|9246_ ;
  assign \new_Sorter100|9347_  = \new_Sorter100|9247_  & \new_Sorter100|9248_ ;
  assign \new_Sorter100|9348_  = \new_Sorter100|9247_  | \new_Sorter100|9248_ ;
  assign \new_Sorter100|9349_  = \new_Sorter100|9249_  & \new_Sorter100|9250_ ;
  assign \new_Sorter100|9350_  = \new_Sorter100|9249_  | \new_Sorter100|9250_ ;
  assign \new_Sorter100|9351_  = \new_Sorter100|9251_  & \new_Sorter100|9252_ ;
  assign \new_Sorter100|9352_  = \new_Sorter100|9251_  | \new_Sorter100|9252_ ;
  assign \new_Sorter100|9353_  = \new_Sorter100|9253_  & \new_Sorter100|9254_ ;
  assign \new_Sorter100|9354_  = \new_Sorter100|9253_  | \new_Sorter100|9254_ ;
  assign \new_Sorter100|9355_  = \new_Sorter100|9255_  & \new_Sorter100|9256_ ;
  assign \new_Sorter100|9356_  = \new_Sorter100|9255_  | \new_Sorter100|9256_ ;
  assign \new_Sorter100|9357_  = \new_Sorter100|9257_  & \new_Sorter100|9258_ ;
  assign \new_Sorter100|9358_  = \new_Sorter100|9257_  | \new_Sorter100|9258_ ;
  assign \new_Sorter100|9359_  = \new_Sorter100|9259_  & \new_Sorter100|9260_ ;
  assign \new_Sorter100|9360_  = \new_Sorter100|9259_  | \new_Sorter100|9260_ ;
  assign \new_Sorter100|9361_  = \new_Sorter100|9261_  & \new_Sorter100|9262_ ;
  assign \new_Sorter100|9362_  = \new_Sorter100|9261_  | \new_Sorter100|9262_ ;
  assign \new_Sorter100|9363_  = \new_Sorter100|9263_  & \new_Sorter100|9264_ ;
  assign \new_Sorter100|9364_  = \new_Sorter100|9263_  | \new_Sorter100|9264_ ;
  assign \new_Sorter100|9365_  = \new_Sorter100|9265_  & \new_Sorter100|9266_ ;
  assign \new_Sorter100|9366_  = \new_Sorter100|9265_  | \new_Sorter100|9266_ ;
  assign \new_Sorter100|9367_  = \new_Sorter100|9267_  & \new_Sorter100|9268_ ;
  assign \new_Sorter100|9368_  = \new_Sorter100|9267_  | \new_Sorter100|9268_ ;
  assign \new_Sorter100|9369_  = \new_Sorter100|9269_  & \new_Sorter100|9270_ ;
  assign \new_Sorter100|9370_  = \new_Sorter100|9269_  | \new_Sorter100|9270_ ;
  assign \new_Sorter100|9371_  = \new_Sorter100|9271_  & \new_Sorter100|9272_ ;
  assign \new_Sorter100|9372_  = \new_Sorter100|9271_  | \new_Sorter100|9272_ ;
  assign \new_Sorter100|9373_  = \new_Sorter100|9273_  & \new_Sorter100|9274_ ;
  assign \new_Sorter100|9374_  = \new_Sorter100|9273_  | \new_Sorter100|9274_ ;
  assign \new_Sorter100|9375_  = \new_Sorter100|9275_  & \new_Sorter100|9276_ ;
  assign \new_Sorter100|9376_  = \new_Sorter100|9275_  | \new_Sorter100|9276_ ;
  assign \new_Sorter100|9377_  = \new_Sorter100|9277_  & \new_Sorter100|9278_ ;
  assign \new_Sorter100|9378_  = \new_Sorter100|9277_  | \new_Sorter100|9278_ ;
  assign \new_Sorter100|9379_  = \new_Sorter100|9279_  & \new_Sorter100|9280_ ;
  assign \new_Sorter100|9380_  = \new_Sorter100|9279_  | \new_Sorter100|9280_ ;
  assign \new_Sorter100|9381_  = \new_Sorter100|9281_  & \new_Sorter100|9282_ ;
  assign \new_Sorter100|9382_  = \new_Sorter100|9281_  | \new_Sorter100|9282_ ;
  assign \new_Sorter100|9383_  = \new_Sorter100|9283_  & \new_Sorter100|9284_ ;
  assign \new_Sorter100|9384_  = \new_Sorter100|9283_  | \new_Sorter100|9284_ ;
  assign \new_Sorter100|9385_  = \new_Sorter100|9285_  & \new_Sorter100|9286_ ;
  assign \new_Sorter100|9386_  = \new_Sorter100|9285_  | \new_Sorter100|9286_ ;
  assign \new_Sorter100|9387_  = \new_Sorter100|9287_  & \new_Sorter100|9288_ ;
  assign \new_Sorter100|9388_  = \new_Sorter100|9287_  | \new_Sorter100|9288_ ;
  assign \new_Sorter100|9389_  = \new_Sorter100|9289_  & \new_Sorter100|9290_ ;
  assign \new_Sorter100|9390_  = \new_Sorter100|9289_  | \new_Sorter100|9290_ ;
  assign \new_Sorter100|9391_  = \new_Sorter100|9291_  & \new_Sorter100|9292_ ;
  assign \new_Sorter100|9392_  = \new_Sorter100|9291_  | \new_Sorter100|9292_ ;
  assign \new_Sorter100|9393_  = \new_Sorter100|9293_  & \new_Sorter100|9294_ ;
  assign \new_Sorter100|9394_  = \new_Sorter100|9293_  | \new_Sorter100|9294_ ;
  assign \new_Sorter100|9395_  = \new_Sorter100|9295_  & \new_Sorter100|9296_ ;
  assign \new_Sorter100|9396_  = \new_Sorter100|9295_  | \new_Sorter100|9296_ ;
  assign \new_Sorter100|9397_  = \new_Sorter100|9297_  & \new_Sorter100|9298_ ;
  assign \new_Sorter100|9398_  = \new_Sorter100|9297_  | \new_Sorter100|9298_ ;
  assign \new_Sorter100|9400_  = \new_Sorter100|9300_  & \new_Sorter100|9301_ ;
  assign \new_Sorter100|9401_  = \new_Sorter100|9300_  | \new_Sorter100|9301_ ;
  assign \new_Sorter100|9402_  = \new_Sorter100|9302_  & \new_Sorter100|9303_ ;
  assign \new_Sorter100|9403_  = \new_Sorter100|9302_  | \new_Sorter100|9303_ ;
  assign \new_Sorter100|9404_  = \new_Sorter100|9304_  & \new_Sorter100|9305_ ;
  assign \new_Sorter100|9405_  = \new_Sorter100|9304_  | \new_Sorter100|9305_ ;
  assign \new_Sorter100|9406_  = \new_Sorter100|9306_  & \new_Sorter100|9307_ ;
  assign \new_Sorter100|9407_  = \new_Sorter100|9306_  | \new_Sorter100|9307_ ;
  assign \new_Sorter100|9408_  = \new_Sorter100|9308_  & \new_Sorter100|9309_ ;
  assign \new_Sorter100|9409_  = \new_Sorter100|9308_  | \new_Sorter100|9309_ ;
  assign \new_Sorter100|9410_  = \new_Sorter100|9310_  & \new_Sorter100|9311_ ;
  assign \new_Sorter100|9411_  = \new_Sorter100|9310_  | \new_Sorter100|9311_ ;
  assign \new_Sorter100|9412_  = \new_Sorter100|9312_  & \new_Sorter100|9313_ ;
  assign \new_Sorter100|9413_  = \new_Sorter100|9312_  | \new_Sorter100|9313_ ;
  assign \new_Sorter100|9414_  = \new_Sorter100|9314_  & \new_Sorter100|9315_ ;
  assign \new_Sorter100|9415_  = \new_Sorter100|9314_  | \new_Sorter100|9315_ ;
  assign \new_Sorter100|9416_  = \new_Sorter100|9316_  & \new_Sorter100|9317_ ;
  assign \new_Sorter100|9417_  = \new_Sorter100|9316_  | \new_Sorter100|9317_ ;
  assign \new_Sorter100|9418_  = \new_Sorter100|9318_  & \new_Sorter100|9319_ ;
  assign \new_Sorter100|9419_  = \new_Sorter100|9318_  | \new_Sorter100|9319_ ;
  assign \new_Sorter100|9420_  = \new_Sorter100|9320_  & \new_Sorter100|9321_ ;
  assign \new_Sorter100|9421_  = \new_Sorter100|9320_  | \new_Sorter100|9321_ ;
  assign \new_Sorter100|9422_  = \new_Sorter100|9322_  & \new_Sorter100|9323_ ;
  assign \new_Sorter100|9423_  = \new_Sorter100|9322_  | \new_Sorter100|9323_ ;
  assign \new_Sorter100|9424_  = \new_Sorter100|9324_  & \new_Sorter100|9325_ ;
  assign \new_Sorter100|9425_  = \new_Sorter100|9324_  | \new_Sorter100|9325_ ;
  assign \new_Sorter100|9426_  = \new_Sorter100|9326_  & \new_Sorter100|9327_ ;
  assign \new_Sorter100|9427_  = \new_Sorter100|9326_  | \new_Sorter100|9327_ ;
  assign \new_Sorter100|9428_  = \new_Sorter100|9328_  & \new_Sorter100|9329_ ;
  assign \new_Sorter100|9429_  = \new_Sorter100|9328_  | \new_Sorter100|9329_ ;
  assign \new_Sorter100|9430_  = \new_Sorter100|9330_  & \new_Sorter100|9331_ ;
  assign \new_Sorter100|9431_  = \new_Sorter100|9330_  | \new_Sorter100|9331_ ;
  assign \new_Sorter100|9432_  = \new_Sorter100|9332_  & \new_Sorter100|9333_ ;
  assign \new_Sorter100|9433_  = \new_Sorter100|9332_  | \new_Sorter100|9333_ ;
  assign \new_Sorter100|9434_  = \new_Sorter100|9334_  & \new_Sorter100|9335_ ;
  assign \new_Sorter100|9435_  = \new_Sorter100|9334_  | \new_Sorter100|9335_ ;
  assign \new_Sorter100|9436_  = \new_Sorter100|9336_  & \new_Sorter100|9337_ ;
  assign \new_Sorter100|9437_  = \new_Sorter100|9336_  | \new_Sorter100|9337_ ;
  assign \new_Sorter100|9438_  = \new_Sorter100|9338_  & \new_Sorter100|9339_ ;
  assign \new_Sorter100|9439_  = \new_Sorter100|9338_  | \new_Sorter100|9339_ ;
  assign \new_Sorter100|9440_  = \new_Sorter100|9340_  & \new_Sorter100|9341_ ;
  assign \new_Sorter100|9441_  = \new_Sorter100|9340_  | \new_Sorter100|9341_ ;
  assign \new_Sorter100|9442_  = \new_Sorter100|9342_  & \new_Sorter100|9343_ ;
  assign \new_Sorter100|9443_  = \new_Sorter100|9342_  | \new_Sorter100|9343_ ;
  assign \new_Sorter100|9444_  = \new_Sorter100|9344_  & \new_Sorter100|9345_ ;
  assign \new_Sorter100|9445_  = \new_Sorter100|9344_  | \new_Sorter100|9345_ ;
  assign \new_Sorter100|9446_  = \new_Sorter100|9346_  & \new_Sorter100|9347_ ;
  assign \new_Sorter100|9447_  = \new_Sorter100|9346_  | \new_Sorter100|9347_ ;
  assign \new_Sorter100|9448_  = \new_Sorter100|9348_  & \new_Sorter100|9349_ ;
  assign \new_Sorter100|9449_  = \new_Sorter100|9348_  | \new_Sorter100|9349_ ;
  assign \new_Sorter100|9450_  = \new_Sorter100|9350_  & \new_Sorter100|9351_ ;
  assign \new_Sorter100|9451_  = \new_Sorter100|9350_  | \new_Sorter100|9351_ ;
  assign \new_Sorter100|9452_  = \new_Sorter100|9352_  & \new_Sorter100|9353_ ;
  assign \new_Sorter100|9453_  = \new_Sorter100|9352_  | \new_Sorter100|9353_ ;
  assign \new_Sorter100|9454_  = \new_Sorter100|9354_  & \new_Sorter100|9355_ ;
  assign \new_Sorter100|9455_  = \new_Sorter100|9354_  | \new_Sorter100|9355_ ;
  assign \new_Sorter100|9456_  = \new_Sorter100|9356_  & \new_Sorter100|9357_ ;
  assign \new_Sorter100|9457_  = \new_Sorter100|9356_  | \new_Sorter100|9357_ ;
  assign \new_Sorter100|9458_  = \new_Sorter100|9358_  & \new_Sorter100|9359_ ;
  assign \new_Sorter100|9459_  = \new_Sorter100|9358_  | \new_Sorter100|9359_ ;
  assign \new_Sorter100|9460_  = \new_Sorter100|9360_  & \new_Sorter100|9361_ ;
  assign \new_Sorter100|9461_  = \new_Sorter100|9360_  | \new_Sorter100|9361_ ;
  assign \new_Sorter100|9462_  = \new_Sorter100|9362_  & \new_Sorter100|9363_ ;
  assign \new_Sorter100|9463_  = \new_Sorter100|9362_  | \new_Sorter100|9363_ ;
  assign \new_Sorter100|9464_  = \new_Sorter100|9364_  & \new_Sorter100|9365_ ;
  assign \new_Sorter100|9465_  = \new_Sorter100|9364_  | \new_Sorter100|9365_ ;
  assign \new_Sorter100|9466_  = \new_Sorter100|9366_  & \new_Sorter100|9367_ ;
  assign \new_Sorter100|9467_  = \new_Sorter100|9366_  | \new_Sorter100|9367_ ;
  assign \new_Sorter100|9468_  = \new_Sorter100|9368_  & \new_Sorter100|9369_ ;
  assign \new_Sorter100|9469_  = \new_Sorter100|9368_  | \new_Sorter100|9369_ ;
  assign \new_Sorter100|9470_  = \new_Sorter100|9370_  & \new_Sorter100|9371_ ;
  assign \new_Sorter100|9471_  = \new_Sorter100|9370_  | \new_Sorter100|9371_ ;
  assign \new_Sorter100|9472_  = \new_Sorter100|9372_  & \new_Sorter100|9373_ ;
  assign \new_Sorter100|9473_  = \new_Sorter100|9372_  | \new_Sorter100|9373_ ;
  assign \new_Sorter100|9474_  = \new_Sorter100|9374_  & \new_Sorter100|9375_ ;
  assign \new_Sorter100|9475_  = \new_Sorter100|9374_  | \new_Sorter100|9375_ ;
  assign \new_Sorter100|9476_  = \new_Sorter100|9376_  & \new_Sorter100|9377_ ;
  assign \new_Sorter100|9477_  = \new_Sorter100|9376_  | \new_Sorter100|9377_ ;
  assign \new_Sorter100|9478_  = \new_Sorter100|9378_  & \new_Sorter100|9379_ ;
  assign \new_Sorter100|9479_  = \new_Sorter100|9378_  | \new_Sorter100|9379_ ;
  assign \new_Sorter100|9480_  = \new_Sorter100|9380_  & \new_Sorter100|9381_ ;
  assign \new_Sorter100|9481_  = \new_Sorter100|9380_  | \new_Sorter100|9381_ ;
  assign \new_Sorter100|9482_  = \new_Sorter100|9382_  & \new_Sorter100|9383_ ;
  assign \new_Sorter100|9483_  = \new_Sorter100|9382_  | \new_Sorter100|9383_ ;
  assign \new_Sorter100|9484_  = \new_Sorter100|9384_  & \new_Sorter100|9385_ ;
  assign \new_Sorter100|9485_  = \new_Sorter100|9384_  | \new_Sorter100|9385_ ;
  assign \new_Sorter100|9486_  = \new_Sorter100|9386_  & \new_Sorter100|9387_ ;
  assign \new_Sorter100|9487_  = \new_Sorter100|9386_  | \new_Sorter100|9387_ ;
  assign \new_Sorter100|9488_  = \new_Sorter100|9388_  & \new_Sorter100|9389_ ;
  assign \new_Sorter100|9489_  = \new_Sorter100|9388_  | \new_Sorter100|9389_ ;
  assign \new_Sorter100|9490_  = \new_Sorter100|9390_  & \new_Sorter100|9391_ ;
  assign \new_Sorter100|9491_  = \new_Sorter100|9390_  | \new_Sorter100|9391_ ;
  assign \new_Sorter100|9492_  = \new_Sorter100|9392_  & \new_Sorter100|9393_ ;
  assign \new_Sorter100|9493_  = \new_Sorter100|9392_  | \new_Sorter100|9393_ ;
  assign \new_Sorter100|9494_  = \new_Sorter100|9394_  & \new_Sorter100|9395_ ;
  assign \new_Sorter100|9495_  = \new_Sorter100|9394_  | \new_Sorter100|9395_ ;
  assign \new_Sorter100|9496_  = \new_Sorter100|9396_  & \new_Sorter100|9397_ ;
  assign \new_Sorter100|9497_  = \new_Sorter100|9396_  | \new_Sorter100|9397_ ;
  assign \new_Sorter100|9498_  = \new_Sorter100|9398_  & \new_Sorter100|9399_ ;
  assign \new_Sorter100|9499_  = \new_Sorter100|9398_  | \new_Sorter100|9399_ ;
  assign \new_Sorter100|9500_  = \new_Sorter100|9400_ ;
  assign \new_Sorter100|9599_  = \new_Sorter100|9499_ ;
  assign \new_Sorter100|9501_  = \new_Sorter100|9401_  & \new_Sorter100|9402_ ;
  assign \new_Sorter100|9502_  = \new_Sorter100|9401_  | \new_Sorter100|9402_ ;
  assign \new_Sorter100|9503_  = \new_Sorter100|9403_  & \new_Sorter100|9404_ ;
  assign \new_Sorter100|9504_  = \new_Sorter100|9403_  | \new_Sorter100|9404_ ;
  assign \new_Sorter100|9505_  = \new_Sorter100|9405_  & \new_Sorter100|9406_ ;
  assign \new_Sorter100|9506_  = \new_Sorter100|9405_  | \new_Sorter100|9406_ ;
  assign \new_Sorter100|9507_  = \new_Sorter100|9407_  & \new_Sorter100|9408_ ;
  assign \new_Sorter100|9508_  = \new_Sorter100|9407_  | \new_Sorter100|9408_ ;
  assign \new_Sorter100|9509_  = \new_Sorter100|9409_  & \new_Sorter100|9410_ ;
  assign \new_Sorter100|9510_  = \new_Sorter100|9409_  | \new_Sorter100|9410_ ;
  assign \new_Sorter100|9511_  = \new_Sorter100|9411_  & \new_Sorter100|9412_ ;
  assign \new_Sorter100|9512_  = \new_Sorter100|9411_  | \new_Sorter100|9412_ ;
  assign \new_Sorter100|9513_  = \new_Sorter100|9413_  & \new_Sorter100|9414_ ;
  assign \new_Sorter100|9514_  = \new_Sorter100|9413_  | \new_Sorter100|9414_ ;
  assign \new_Sorter100|9515_  = \new_Sorter100|9415_  & \new_Sorter100|9416_ ;
  assign \new_Sorter100|9516_  = \new_Sorter100|9415_  | \new_Sorter100|9416_ ;
  assign \new_Sorter100|9517_  = \new_Sorter100|9417_  & \new_Sorter100|9418_ ;
  assign \new_Sorter100|9518_  = \new_Sorter100|9417_  | \new_Sorter100|9418_ ;
  assign \new_Sorter100|9519_  = \new_Sorter100|9419_  & \new_Sorter100|9420_ ;
  assign \new_Sorter100|9520_  = \new_Sorter100|9419_  | \new_Sorter100|9420_ ;
  assign \new_Sorter100|9521_  = \new_Sorter100|9421_  & \new_Sorter100|9422_ ;
  assign \new_Sorter100|9522_  = \new_Sorter100|9421_  | \new_Sorter100|9422_ ;
  assign \new_Sorter100|9523_  = \new_Sorter100|9423_  & \new_Sorter100|9424_ ;
  assign \new_Sorter100|9524_  = \new_Sorter100|9423_  | \new_Sorter100|9424_ ;
  assign \new_Sorter100|9525_  = \new_Sorter100|9425_  & \new_Sorter100|9426_ ;
  assign \new_Sorter100|9526_  = \new_Sorter100|9425_  | \new_Sorter100|9426_ ;
  assign \new_Sorter100|9527_  = \new_Sorter100|9427_  & \new_Sorter100|9428_ ;
  assign \new_Sorter100|9528_  = \new_Sorter100|9427_  | \new_Sorter100|9428_ ;
  assign \new_Sorter100|9529_  = \new_Sorter100|9429_  & \new_Sorter100|9430_ ;
  assign \new_Sorter100|9530_  = \new_Sorter100|9429_  | \new_Sorter100|9430_ ;
  assign \new_Sorter100|9531_  = \new_Sorter100|9431_  & \new_Sorter100|9432_ ;
  assign \new_Sorter100|9532_  = \new_Sorter100|9431_  | \new_Sorter100|9432_ ;
  assign \new_Sorter100|9533_  = \new_Sorter100|9433_  & \new_Sorter100|9434_ ;
  assign \new_Sorter100|9534_  = \new_Sorter100|9433_  | \new_Sorter100|9434_ ;
  assign \new_Sorter100|9535_  = \new_Sorter100|9435_  & \new_Sorter100|9436_ ;
  assign \new_Sorter100|9536_  = \new_Sorter100|9435_  | \new_Sorter100|9436_ ;
  assign \new_Sorter100|9537_  = \new_Sorter100|9437_  & \new_Sorter100|9438_ ;
  assign \new_Sorter100|9538_  = \new_Sorter100|9437_  | \new_Sorter100|9438_ ;
  assign \new_Sorter100|9539_  = \new_Sorter100|9439_  & \new_Sorter100|9440_ ;
  assign \new_Sorter100|9540_  = \new_Sorter100|9439_  | \new_Sorter100|9440_ ;
  assign \new_Sorter100|9541_  = \new_Sorter100|9441_  & \new_Sorter100|9442_ ;
  assign \new_Sorter100|9542_  = \new_Sorter100|9441_  | \new_Sorter100|9442_ ;
  assign \new_Sorter100|9543_  = \new_Sorter100|9443_  & \new_Sorter100|9444_ ;
  assign \new_Sorter100|9544_  = \new_Sorter100|9443_  | \new_Sorter100|9444_ ;
  assign \new_Sorter100|9545_  = \new_Sorter100|9445_  & \new_Sorter100|9446_ ;
  assign \new_Sorter100|9546_  = \new_Sorter100|9445_  | \new_Sorter100|9446_ ;
  assign \new_Sorter100|9547_  = \new_Sorter100|9447_  & \new_Sorter100|9448_ ;
  assign \new_Sorter100|9548_  = \new_Sorter100|9447_  | \new_Sorter100|9448_ ;
  assign \new_Sorter100|9549_  = \new_Sorter100|9449_  & \new_Sorter100|9450_ ;
  assign \new_Sorter100|9550_  = \new_Sorter100|9449_  | \new_Sorter100|9450_ ;
  assign \new_Sorter100|9551_  = \new_Sorter100|9451_  & \new_Sorter100|9452_ ;
  assign \new_Sorter100|9552_  = \new_Sorter100|9451_  | \new_Sorter100|9452_ ;
  assign \new_Sorter100|9553_  = \new_Sorter100|9453_  & \new_Sorter100|9454_ ;
  assign \new_Sorter100|9554_  = \new_Sorter100|9453_  | \new_Sorter100|9454_ ;
  assign \new_Sorter100|9555_  = \new_Sorter100|9455_  & \new_Sorter100|9456_ ;
  assign \new_Sorter100|9556_  = \new_Sorter100|9455_  | \new_Sorter100|9456_ ;
  assign \new_Sorter100|9557_  = \new_Sorter100|9457_  & \new_Sorter100|9458_ ;
  assign \new_Sorter100|9558_  = \new_Sorter100|9457_  | \new_Sorter100|9458_ ;
  assign \new_Sorter100|9559_  = \new_Sorter100|9459_  & \new_Sorter100|9460_ ;
  assign \new_Sorter100|9560_  = \new_Sorter100|9459_  | \new_Sorter100|9460_ ;
  assign \new_Sorter100|9561_  = \new_Sorter100|9461_  & \new_Sorter100|9462_ ;
  assign \new_Sorter100|9562_  = \new_Sorter100|9461_  | \new_Sorter100|9462_ ;
  assign \new_Sorter100|9563_  = \new_Sorter100|9463_  & \new_Sorter100|9464_ ;
  assign \new_Sorter100|9564_  = \new_Sorter100|9463_  | \new_Sorter100|9464_ ;
  assign \new_Sorter100|9565_  = \new_Sorter100|9465_  & \new_Sorter100|9466_ ;
  assign \new_Sorter100|9566_  = \new_Sorter100|9465_  | \new_Sorter100|9466_ ;
  assign \new_Sorter100|9567_  = \new_Sorter100|9467_  & \new_Sorter100|9468_ ;
  assign \new_Sorter100|9568_  = \new_Sorter100|9467_  | \new_Sorter100|9468_ ;
  assign \new_Sorter100|9569_  = \new_Sorter100|9469_  & \new_Sorter100|9470_ ;
  assign \new_Sorter100|9570_  = \new_Sorter100|9469_  | \new_Sorter100|9470_ ;
  assign \new_Sorter100|9571_  = \new_Sorter100|9471_  & \new_Sorter100|9472_ ;
  assign \new_Sorter100|9572_  = \new_Sorter100|9471_  | \new_Sorter100|9472_ ;
  assign \new_Sorter100|9573_  = \new_Sorter100|9473_  & \new_Sorter100|9474_ ;
  assign \new_Sorter100|9574_  = \new_Sorter100|9473_  | \new_Sorter100|9474_ ;
  assign \new_Sorter100|9575_  = \new_Sorter100|9475_  & \new_Sorter100|9476_ ;
  assign \new_Sorter100|9576_  = \new_Sorter100|9475_  | \new_Sorter100|9476_ ;
  assign \new_Sorter100|9577_  = \new_Sorter100|9477_  & \new_Sorter100|9478_ ;
  assign \new_Sorter100|9578_  = \new_Sorter100|9477_  | \new_Sorter100|9478_ ;
  assign \new_Sorter100|9579_  = \new_Sorter100|9479_  & \new_Sorter100|9480_ ;
  assign \new_Sorter100|9580_  = \new_Sorter100|9479_  | \new_Sorter100|9480_ ;
  assign \new_Sorter100|9581_  = \new_Sorter100|9481_  & \new_Sorter100|9482_ ;
  assign \new_Sorter100|9582_  = \new_Sorter100|9481_  | \new_Sorter100|9482_ ;
  assign \new_Sorter100|9583_  = \new_Sorter100|9483_  & \new_Sorter100|9484_ ;
  assign \new_Sorter100|9584_  = \new_Sorter100|9483_  | \new_Sorter100|9484_ ;
  assign \new_Sorter100|9585_  = \new_Sorter100|9485_  & \new_Sorter100|9486_ ;
  assign \new_Sorter100|9586_  = \new_Sorter100|9485_  | \new_Sorter100|9486_ ;
  assign \new_Sorter100|9587_  = \new_Sorter100|9487_  & \new_Sorter100|9488_ ;
  assign \new_Sorter100|9588_  = \new_Sorter100|9487_  | \new_Sorter100|9488_ ;
  assign \new_Sorter100|9589_  = \new_Sorter100|9489_  & \new_Sorter100|9490_ ;
  assign \new_Sorter100|9590_  = \new_Sorter100|9489_  | \new_Sorter100|9490_ ;
  assign \new_Sorter100|9591_  = \new_Sorter100|9491_  & \new_Sorter100|9492_ ;
  assign \new_Sorter100|9592_  = \new_Sorter100|9491_  | \new_Sorter100|9492_ ;
  assign \new_Sorter100|9593_  = \new_Sorter100|9493_  & \new_Sorter100|9494_ ;
  assign \new_Sorter100|9594_  = \new_Sorter100|9493_  | \new_Sorter100|9494_ ;
  assign \new_Sorter100|9595_  = \new_Sorter100|9495_  & \new_Sorter100|9496_ ;
  assign \new_Sorter100|9596_  = \new_Sorter100|9495_  | \new_Sorter100|9496_ ;
  assign \new_Sorter100|9597_  = \new_Sorter100|9497_  & \new_Sorter100|9498_ ;
  assign \new_Sorter100|9598_  = \new_Sorter100|9497_  | \new_Sorter100|9498_ ;
  assign \new_Sorter100|9600_  = \new_Sorter100|9500_  & \new_Sorter100|9501_ ;
  assign \new_Sorter100|9601_  = \new_Sorter100|9500_  | \new_Sorter100|9501_ ;
  assign \new_Sorter100|9602_  = \new_Sorter100|9502_  & \new_Sorter100|9503_ ;
  assign \new_Sorter100|9603_  = \new_Sorter100|9502_  | \new_Sorter100|9503_ ;
  assign \new_Sorter100|9604_  = \new_Sorter100|9504_  & \new_Sorter100|9505_ ;
  assign \new_Sorter100|9605_  = \new_Sorter100|9504_  | \new_Sorter100|9505_ ;
  assign \new_Sorter100|9606_  = \new_Sorter100|9506_  & \new_Sorter100|9507_ ;
  assign \new_Sorter100|9607_  = \new_Sorter100|9506_  | \new_Sorter100|9507_ ;
  assign \new_Sorter100|9608_  = \new_Sorter100|9508_  & \new_Sorter100|9509_ ;
  assign \new_Sorter100|9609_  = \new_Sorter100|9508_  | \new_Sorter100|9509_ ;
  assign \new_Sorter100|9610_  = \new_Sorter100|9510_  & \new_Sorter100|9511_ ;
  assign \new_Sorter100|9611_  = \new_Sorter100|9510_  | \new_Sorter100|9511_ ;
  assign \new_Sorter100|9612_  = \new_Sorter100|9512_  & \new_Sorter100|9513_ ;
  assign \new_Sorter100|9613_  = \new_Sorter100|9512_  | \new_Sorter100|9513_ ;
  assign \new_Sorter100|9614_  = \new_Sorter100|9514_  & \new_Sorter100|9515_ ;
  assign \new_Sorter100|9615_  = \new_Sorter100|9514_  | \new_Sorter100|9515_ ;
  assign \new_Sorter100|9616_  = \new_Sorter100|9516_  & \new_Sorter100|9517_ ;
  assign \new_Sorter100|9617_  = \new_Sorter100|9516_  | \new_Sorter100|9517_ ;
  assign \new_Sorter100|9618_  = \new_Sorter100|9518_  & \new_Sorter100|9519_ ;
  assign \new_Sorter100|9619_  = \new_Sorter100|9518_  | \new_Sorter100|9519_ ;
  assign \new_Sorter100|9620_  = \new_Sorter100|9520_  & \new_Sorter100|9521_ ;
  assign \new_Sorter100|9621_  = \new_Sorter100|9520_  | \new_Sorter100|9521_ ;
  assign \new_Sorter100|9622_  = \new_Sorter100|9522_  & \new_Sorter100|9523_ ;
  assign \new_Sorter100|9623_  = \new_Sorter100|9522_  | \new_Sorter100|9523_ ;
  assign \new_Sorter100|9624_  = \new_Sorter100|9524_  & \new_Sorter100|9525_ ;
  assign \new_Sorter100|9625_  = \new_Sorter100|9524_  | \new_Sorter100|9525_ ;
  assign \new_Sorter100|9626_  = \new_Sorter100|9526_  & \new_Sorter100|9527_ ;
  assign \new_Sorter100|9627_  = \new_Sorter100|9526_  | \new_Sorter100|9527_ ;
  assign \new_Sorter100|9628_  = \new_Sorter100|9528_  & \new_Sorter100|9529_ ;
  assign \new_Sorter100|9629_  = \new_Sorter100|9528_  | \new_Sorter100|9529_ ;
  assign \new_Sorter100|9630_  = \new_Sorter100|9530_  & \new_Sorter100|9531_ ;
  assign \new_Sorter100|9631_  = \new_Sorter100|9530_  | \new_Sorter100|9531_ ;
  assign \new_Sorter100|9632_  = \new_Sorter100|9532_  & \new_Sorter100|9533_ ;
  assign \new_Sorter100|9633_  = \new_Sorter100|9532_  | \new_Sorter100|9533_ ;
  assign \new_Sorter100|9634_  = \new_Sorter100|9534_  & \new_Sorter100|9535_ ;
  assign \new_Sorter100|9635_  = \new_Sorter100|9534_  | \new_Sorter100|9535_ ;
  assign \new_Sorter100|9636_  = \new_Sorter100|9536_  & \new_Sorter100|9537_ ;
  assign \new_Sorter100|9637_  = \new_Sorter100|9536_  | \new_Sorter100|9537_ ;
  assign \new_Sorter100|9638_  = \new_Sorter100|9538_  & \new_Sorter100|9539_ ;
  assign \new_Sorter100|9639_  = \new_Sorter100|9538_  | \new_Sorter100|9539_ ;
  assign \new_Sorter100|9640_  = \new_Sorter100|9540_  & \new_Sorter100|9541_ ;
  assign \new_Sorter100|9641_  = \new_Sorter100|9540_  | \new_Sorter100|9541_ ;
  assign \new_Sorter100|9642_  = \new_Sorter100|9542_  & \new_Sorter100|9543_ ;
  assign \new_Sorter100|9643_  = \new_Sorter100|9542_  | \new_Sorter100|9543_ ;
  assign \new_Sorter100|9644_  = \new_Sorter100|9544_  & \new_Sorter100|9545_ ;
  assign \new_Sorter100|9645_  = \new_Sorter100|9544_  | \new_Sorter100|9545_ ;
  assign \new_Sorter100|9646_  = \new_Sorter100|9546_  & \new_Sorter100|9547_ ;
  assign \new_Sorter100|9647_  = \new_Sorter100|9546_  | \new_Sorter100|9547_ ;
  assign \new_Sorter100|9648_  = \new_Sorter100|9548_  & \new_Sorter100|9549_ ;
  assign \new_Sorter100|9649_  = \new_Sorter100|9548_  | \new_Sorter100|9549_ ;
  assign \new_Sorter100|9650_  = \new_Sorter100|9550_  & \new_Sorter100|9551_ ;
  assign \new_Sorter100|9651_  = \new_Sorter100|9550_  | \new_Sorter100|9551_ ;
  assign \new_Sorter100|9652_  = \new_Sorter100|9552_  & \new_Sorter100|9553_ ;
  assign \new_Sorter100|9653_  = \new_Sorter100|9552_  | \new_Sorter100|9553_ ;
  assign \new_Sorter100|9654_  = \new_Sorter100|9554_  & \new_Sorter100|9555_ ;
  assign \new_Sorter100|9655_  = \new_Sorter100|9554_  | \new_Sorter100|9555_ ;
  assign \new_Sorter100|9656_  = \new_Sorter100|9556_  & \new_Sorter100|9557_ ;
  assign \new_Sorter100|9657_  = \new_Sorter100|9556_  | \new_Sorter100|9557_ ;
  assign \new_Sorter100|9658_  = \new_Sorter100|9558_  & \new_Sorter100|9559_ ;
  assign \new_Sorter100|9659_  = \new_Sorter100|9558_  | \new_Sorter100|9559_ ;
  assign \new_Sorter100|9660_  = \new_Sorter100|9560_  & \new_Sorter100|9561_ ;
  assign \new_Sorter100|9661_  = \new_Sorter100|9560_  | \new_Sorter100|9561_ ;
  assign \new_Sorter100|9662_  = \new_Sorter100|9562_  & \new_Sorter100|9563_ ;
  assign \new_Sorter100|9663_  = \new_Sorter100|9562_  | \new_Sorter100|9563_ ;
  assign \new_Sorter100|9664_  = \new_Sorter100|9564_  & \new_Sorter100|9565_ ;
  assign \new_Sorter100|9665_  = \new_Sorter100|9564_  | \new_Sorter100|9565_ ;
  assign \new_Sorter100|9666_  = \new_Sorter100|9566_  & \new_Sorter100|9567_ ;
  assign \new_Sorter100|9667_  = \new_Sorter100|9566_  | \new_Sorter100|9567_ ;
  assign \new_Sorter100|9668_  = \new_Sorter100|9568_  & \new_Sorter100|9569_ ;
  assign \new_Sorter100|9669_  = \new_Sorter100|9568_  | \new_Sorter100|9569_ ;
  assign \new_Sorter100|9670_  = \new_Sorter100|9570_  & \new_Sorter100|9571_ ;
  assign \new_Sorter100|9671_  = \new_Sorter100|9570_  | \new_Sorter100|9571_ ;
  assign \new_Sorter100|9672_  = \new_Sorter100|9572_  & \new_Sorter100|9573_ ;
  assign \new_Sorter100|9673_  = \new_Sorter100|9572_  | \new_Sorter100|9573_ ;
  assign \new_Sorter100|9674_  = \new_Sorter100|9574_  & \new_Sorter100|9575_ ;
  assign \new_Sorter100|9675_  = \new_Sorter100|9574_  | \new_Sorter100|9575_ ;
  assign \new_Sorter100|9676_  = \new_Sorter100|9576_  & \new_Sorter100|9577_ ;
  assign \new_Sorter100|9677_  = \new_Sorter100|9576_  | \new_Sorter100|9577_ ;
  assign \new_Sorter100|9678_  = \new_Sorter100|9578_  & \new_Sorter100|9579_ ;
  assign \new_Sorter100|9679_  = \new_Sorter100|9578_  | \new_Sorter100|9579_ ;
  assign \new_Sorter100|9680_  = \new_Sorter100|9580_  & \new_Sorter100|9581_ ;
  assign \new_Sorter100|9681_  = \new_Sorter100|9580_  | \new_Sorter100|9581_ ;
  assign \new_Sorter100|9682_  = \new_Sorter100|9582_  & \new_Sorter100|9583_ ;
  assign \new_Sorter100|9683_  = \new_Sorter100|9582_  | \new_Sorter100|9583_ ;
  assign \new_Sorter100|9684_  = \new_Sorter100|9584_  & \new_Sorter100|9585_ ;
  assign \new_Sorter100|9685_  = \new_Sorter100|9584_  | \new_Sorter100|9585_ ;
  assign \new_Sorter100|9686_  = \new_Sorter100|9586_  & \new_Sorter100|9587_ ;
  assign \new_Sorter100|9687_  = \new_Sorter100|9586_  | \new_Sorter100|9587_ ;
  assign \new_Sorter100|9688_  = \new_Sorter100|9588_  & \new_Sorter100|9589_ ;
  assign \new_Sorter100|9689_  = \new_Sorter100|9588_  | \new_Sorter100|9589_ ;
  assign \new_Sorter100|9690_  = \new_Sorter100|9590_  & \new_Sorter100|9591_ ;
  assign \new_Sorter100|9691_  = \new_Sorter100|9590_  | \new_Sorter100|9591_ ;
  assign \new_Sorter100|9692_  = \new_Sorter100|9592_  & \new_Sorter100|9593_ ;
  assign \new_Sorter100|9693_  = \new_Sorter100|9592_  | \new_Sorter100|9593_ ;
  assign \new_Sorter100|9694_  = \new_Sorter100|9594_  & \new_Sorter100|9595_ ;
  assign \new_Sorter100|9695_  = \new_Sorter100|9594_  | \new_Sorter100|9595_ ;
  assign \new_Sorter100|9696_  = \new_Sorter100|9596_  & \new_Sorter100|9597_ ;
  assign \new_Sorter100|9697_  = \new_Sorter100|9596_  | \new_Sorter100|9597_ ;
  assign \new_Sorter100|9698_  = \new_Sorter100|9598_  & \new_Sorter100|9599_ ;
  assign \new_Sorter100|9699_  = \new_Sorter100|9598_  | \new_Sorter100|9599_ ;
  assign \new_Sorter100|9700_  = \new_Sorter100|9600_ ;
  assign \new_Sorter100|9799_  = \new_Sorter100|9699_ ;
  assign \new_Sorter100|9701_  = \new_Sorter100|9601_  & \new_Sorter100|9602_ ;
  assign \new_Sorter100|9702_  = \new_Sorter100|9601_  | \new_Sorter100|9602_ ;
  assign \new_Sorter100|9703_  = \new_Sorter100|9603_  & \new_Sorter100|9604_ ;
  assign \new_Sorter100|9704_  = \new_Sorter100|9603_  | \new_Sorter100|9604_ ;
  assign \new_Sorter100|9705_  = \new_Sorter100|9605_  & \new_Sorter100|9606_ ;
  assign \new_Sorter100|9706_  = \new_Sorter100|9605_  | \new_Sorter100|9606_ ;
  assign \new_Sorter100|9707_  = \new_Sorter100|9607_  & \new_Sorter100|9608_ ;
  assign \new_Sorter100|9708_  = \new_Sorter100|9607_  | \new_Sorter100|9608_ ;
  assign \new_Sorter100|9709_  = \new_Sorter100|9609_  & \new_Sorter100|9610_ ;
  assign \new_Sorter100|9710_  = \new_Sorter100|9609_  | \new_Sorter100|9610_ ;
  assign \new_Sorter100|9711_  = \new_Sorter100|9611_  & \new_Sorter100|9612_ ;
  assign \new_Sorter100|9712_  = \new_Sorter100|9611_  | \new_Sorter100|9612_ ;
  assign \new_Sorter100|9713_  = \new_Sorter100|9613_  & \new_Sorter100|9614_ ;
  assign \new_Sorter100|9714_  = \new_Sorter100|9613_  | \new_Sorter100|9614_ ;
  assign \new_Sorter100|9715_  = \new_Sorter100|9615_  & \new_Sorter100|9616_ ;
  assign \new_Sorter100|9716_  = \new_Sorter100|9615_  | \new_Sorter100|9616_ ;
  assign \new_Sorter100|9717_  = \new_Sorter100|9617_  & \new_Sorter100|9618_ ;
  assign \new_Sorter100|9718_  = \new_Sorter100|9617_  | \new_Sorter100|9618_ ;
  assign \new_Sorter100|9719_  = \new_Sorter100|9619_  & \new_Sorter100|9620_ ;
  assign \new_Sorter100|9720_  = \new_Sorter100|9619_  | \new_Sorter100|9620_ ;
  assign \new_Sorter100|9721_  = \new_Sorter100|9621_  & \new_Sorter100|9622_ ;
  assign \new_Sorter100|9722_  = \new_Sorter100|9621_  | \new_Sorter100|9622_ ;
  assign \new_Sorter100|9723_  = \new_Sorter100|9623_  & \new_Sorter100|9624_ ;
  assign \new_Sorter100|9724_  = \new_Sorter100|9623_  | \new_Sorter100|9624_ ;
  assign \new_Sorter100|9725_  = \new_Sorter100|9625_  & \new_Sorter100|9626_ ;
  assign \new_Sorter100|9726_  = \new_Sorter100|9625_  | \new_Sorter100|9626_ ;
  assign \new_Sorter100|9727_  = \new_Sorter100|9627_  & \new_Sorter100|9628_ ;
  assign \new_Sorter100|9728_  = \new_Sorter100|9627_  | \new_Sorter100|9628_ ;
  assign \new_Sorter100|9729_  = \new_Sorter100|9629_  & \new_Sorter100|9630_ ;
  assign \new_Sorter100|9730_  = \new_Sorter100|9629_  | \new_Sorter100|9630_ ;
  assign \new_Sorter100|9731_  = \new_Sorter100|9631_  & \new_Sorter100|9632_ ;
  assign \new_Sorter100|9732_  = \new_Sorter100|9631_  | \new_Sorter100|9632_ ;
  assign \new_Sorter100|9733_  = \new_Sorter100|9633_  & \new_Sorter100|9634_ ;
  assign \new_Sorter100|9734_  = \new_Sorter100|9633_  | \new_Sorter100|9634_ ;
  assign \new_Sorter100|9735_  = \new_Sorter100|9635_  & \new_Sorter100|9636_ ;
  assign \new_Sorter100|9736_  = \new_Sorter100|9635_  | \new_Sorter100|9636_ ;
  assign \new_Sorter100|9737_  = \new_Sorter100|9637_  & \new_Sorter100|9638_ ;
  assign \new_Sorter100|9738_  = \new_Sorter100|9637_  | \new_Sorter100|9638_ ;
  assign \new_Sorter100|9739_  = \new_Sorter100|9639_  & \new_Sorter100|9640_ ;
  assign \new_Sorter100|9740_  = \new_Sorter100|9639_  | \new_Sorter100|9640_ ;
  assign \new_Sorter100|9741_  = \new_Sorter100|9641_  & \new_Sorter100|9642_ ;
  assign \new_Sorter100|9742_  = \new_Sorter100|9641_  | \new_Sorter100|9642_ ;
  assign \new_Sorter100|9743_  = \new_Sorter100|9643_  & \new_Sorter100|9644_ ;
  assign \new_Sorter100|9744_  = \new_Sorter100|9643_  | \new_Sorter100|9644_ ;
  assign \new_Sorter100|9745_  = \new_Sorter100|9645_  & \new_Sorter100|9646_ ;
  assign \new_Sorter100|9746_  = \new_Sorter100|9645_  | \new_Sorter100|9646_ ;
  assign \new_Sorter100|9747_  = \new_Sorter100|9647_  & \new_Sorter100|9648_ ;
  assign \new_Sorter100|9748_  = \new_Sorter100|9647_  | \new_Sorter100|9648_ ;
  assign \new_Sorter100|9749_  = \new_Sorter100|9649_  & \new_Sorter100|9650_ ;
  assign \new_Sorter100|9750_  = \new_Sorter100|9649_  | \new_Sorter100|9650_ ;
  assign \new_Sorter100|9751_  = \new_Sorter100|9651_  & \new_Sorter100|9652_ ;
  assign \new_Sorter100|9752_  = \new_Sorter100|9651_  | \new_Sorter100|9652_ ;
  assign \new_Sorter100|9753_  = \new_Sorter100|9653_  & \new_Sorter100|9654_ ;
  assign \new_Sorter100|9754_  = \new_Sorter100|9653_  | \new_Sorter100|9654_ ;
  assign \new_Sorter100|9755_  = \new_Sorter100|9655_  & \new_Sorter100|9656_ ;
  assign \new_Sorter100|9756_  = \new_Sorter100|9655_  | \new_Sorter100|9656_ ;
  assign \new_Sorter100|9757_  = \new_Sorter100|9657_  & \new_Sorter100|9658_ ;
  assign \new_Sorter100|9758_  = \new_Sorter100|9657_  | \new_Sorter100|9658_ ;
  assign \new_Sorter100|9759_  = \new_Sorter100|9659_  & \new_Sorter100|9660_ ;
  assign \new_Sorter100|9760_  = \new_Sorter100|9659_  | \new_Sorter100|9660_ ;
  assign \new_Sorter100|9761_  = \new_Sorter100|9661_  & \new_Sorter100|9662_ ;
  assign \new_Sorter100|9762_  = \new_Sorter100|9661_  | \new_Sorter100|9662_ ;
  assign \new_Sorter100|9763_  = \new_Sorter100|9663_  & \new_Sorter100|9664_ ;
  assign \new_Sorter100|9764_  = \new_Sorter100|9663_  | \new_Sorter100|9664_ ;
  assign \new_Sorter100|9765_  = \new_Sorter100|9665_  & \new_Sorter100|9666_ ;
  assign \new_Sorter100|9766_  = \new_Sorter100|9665_  | \new_Sorter100|9666_ ;
  assign \new_Sorter100|9767_  = \new_Sorter100|9667_  & \new_Sorter100|9668_ ;
  assign \new_Sorter100|9768_  = \new_Sorter100|9667_  | \new_Sorter100|9668_ ;
  assign \new_Sorter100|9769_  = \new_Sorter100|9669_  & \new_Sorter100|9670_ ;
  assign \new_Sorter100|9770_  = \new_Sorter100|9669_  | \new_Sorter100|9670_ ;
  assign \new_Sorter100|9771_  = \new_Sorter100|9671_  & \new_Sorter100|9672_ ;
  assign \new_Sorter100|9772_  = \new_Sorter100|9671_  | \new_Sorter100|9672_ ;
  assign \new_Sorter100|9773_  = \new_Sorter100|9673_  & \new_Sorter100|9674_ ;
  assign \new_Sorter100|9774_  = \new_Sorter100|9673_  | \new_Sorter100|9674_ ;
  assign \new_Sorter100|9775_  = \new_Sorter100|9675_  & \new_Sorter100|9676_ ;
  assign \new_Sorter100|9776_  = \new_Sorter100|9675_  | \new_Sorter100|9676_ ;
  assign \new_Sorter100|9777_  = \new_Sorter100|9677_  & \new_Sorter100|9678_ ;
  assign \new_Sorter100|9778_  = \new_Sorter100|9677_  | \new_Sorter100|9678_ ;
  assign \new_Sorter100|9779_  = \new_Sorter100|9679_  & \new_Sorter100|9680_ ;
  assign \new_Sorter100|9780_  = \new_Sorter100|9679_  | \new_Sorter100|9680_ ;
  assign \new_Sorter100|9781_  = \new_Sorter100|9681_  & \new_Sorter100|9682_ ;
  assign \new_Sorter100|9782_  = \new_Sorter100|9681_  | \new_Sorter100|9682_ ;
  assign \new_Sorter100|9783_  = \new_Sorter100|9683_  & \new_Sorter100|9684_ ;
  assign \new_Sorter100|9784_  = \new_Sorter100|9683_  | \new_Sorter100|9684_ ;
  assign \new_Sorter100|9785_  = \new_Sorter100|9685_  & \new_Sorter100|9686_ ;
  assign \new_Sorter100|9786_  = \new_Sorter100|9685_  | \new_Sorter100|9686_ ;
  assign \new_Sorter100|9787_  = \new_Sorter100|9687_  & \new_Sorter100|9688_ ;
  assign \new_Sorter100|9788_  = \new_Sorter100|9687_  | \new_Sorter100|9688_ ;
  assign \new_Sorter100|9789_  = \new_Sorter100|9689_  & \new_Sorter100|9690_ ;
  assign \new_Sorter100|9790_  = \new_Sorter100|9689_  | \new_Sorter100|9690_ ;
  assign \new_Sorter100|9791_  = \new_Sorter100|9691_  & \new_Sorter100|9692_ ;
  assign \new_Sorter100|9792_  = \new_Sorter100|9691_  | \new_Sorter100|9692_ ;
  assign \new_Sorter100|9793_  = \new_Sorter100|9693_  & \new_Sorter100|9694_ ;
  assign \new_Sorter100|9794_  = \new_Sorter100|9693_  | \new_Sorter100|9694_ ;
  assign \new_Sorter100|9795_  = \new_Sorter100|9695_  & \new_Sorter100|9696_ ;
  assign \new_Sorter100|9796_  = \new_Sorter100|9695_  | \new_Sorter100|9696_ ;
  assign \new_Sorter100|9797_  = \new_Sorter100|9697_  & \new_Sorter100|9698_ ;
  assign \new_Sorter100|9798_  = \new_Sorter100|9697_  | \new_Sorter100|9698_ ;
  assign \new_Sorter100|9800_  = \new_Sorter100|9700_  & \new_Sorter100|9701_ ;
  assign \new_Sorter100|9801_  = \new_Sorter100|9700_  | \new_Sorter100|9701_ ;
  assign \new_Sorter100|9802_  = \new_Sorter100|9702_  & \new_Sorter100|9703_ ;
  assign \new_Sorter100|9803_  = \new_Sorter100|9702_  | \new_Sorter100|9703_ ;
  assign \new_Sorter100|9804_  = \new_Sorter100|9704_  & \new_Sorter100|9705_ ;
  assign \new_Sorter100|9805_  = \new_Sorter100|9704_  | \new_Sorter100|9705_ ;
  assign \new_Sorter100|9806_  = \new_Sorter100|9706_  & \new_Sorter100|9707_ ;
  assign \new_Sorter100|9807_  = \new_Sorter100|9706_  | \new_Sorter100|9707_ ;
  assign \new_Sorter100|9808_  = \new_Sorter100|9708_  & \new_Sorter100|9709_ ;
  assign \new_Sorter100|9809_  = \new_Sorter100|9708_  | \new_Sorter100|9709_ ;
  assign \new_Sorter100|9810_  = \new_Sorter100|9710_  & \new_Sorter100|9711_ ;
  assign \new_Sorter100|9811_  = \new_Sorter100|9710_  | \new_Sorter100|9711_ ;
  assign \new_Sorter100|9812_  = \new_Sorter100|9712_  & \new_Sorter100|9713_ ;
  assign \new_Sorter100|9813_  = \new_Sorter100|9712_  | \new_Sorter100|9713_ ;
  assign \new_Sorter100|9814_  = \new_Sorter100|9714_  & \new_Sorter100|9715_ ;
  assign \new_Sorter100|9815_  = \new_Sorter100|9714_  | \new_Sorter100|9715_ ;
  assign \new_Sorter100|9816_  = \new_Sorter100|9716_  & \new_Sorter100|9717_ ;
  assign \new_Sorter100|9817_  = \new_Sorter100|9716_  | \new_Sorter100|9717_ ;
  assign \new_Sorter100|9818_  = \new_Sorter100|9718_  & \new_Sorter100|9719_ ;
  assign \new_Sorter100|9819_  = \new_Sorter100|9718_  | \new_Sorter100|9719_ ;
  assign \new_Sorter100|9820_  = \new_Sorter100|9720_  & \new_Sorter100|9721_ ;
  assign \new_Sorter100|9821_  = \new_Sorter100|9720_  | \new_Sorter100|9721_ ;
  assign \new_Sorter100|9822_  = \new_Sorter100|9722_  & \new_Sorter100|9723_ ;
  assign \new_Sorter100|9823_  = \new_Sorter100|9722_  | \new_Sorter100|9723_ ;
  assign \new_Sorter100|9824_  = \new_Sorter100|9724_  & \new_Sorter100|9725_ ;
  assign \new_Sorter100|9825_  = \new_Sorter100|9724_  | \new_Sorter100|9725_ ;
  assign \new_Sorter100|9826_  = \new_Sorter100|9726_  & \new_Sorter100|9727_ ;
  assign \new_Sorter100|9827_  = \new_Sorter100|9726_  | \new_Sorter100|9727_ ;
  assign \new_Sorter100|9828_  = \new_Sorter100|9728_  & \new_Sorter100|9729_ ;
  assign \new_Sorter100|9829_  = \new_Sorter100|9728_  | \new_Sorter100|9729_ ;
  assign \new_Sorter100|9830_  = \new_Sorter100|9730_  & \new_Sorter100|9731_ ;
  assign \new_Sorter100|9831_  = \new_Sorter100|9730_  | \new_Sorter100|9731_ ;
  assign \new_Sorter100|9832_  = \new_Sorter100|9732_  & \new_Sorter100|9733_ ;
  assign \new_Sorter100|9833_  = \new_Sorter100|9732_  | \new_Sorter100|9733_ ;
  assign \new_Sorter100|9834_  = \new_Sorter100|9734_  & \new_Sorter100|9735_ ;
  assign \new_Sorter100|9835_  = \new_Sorter100|9734_  | \new_Sorter100|9735_ ;
  assign \new_Sorter100|9836_  = \new_Sorter100|9736_  & \new_Sorter100|9737_ ;
  assign \new_Sorter100|9837_  = \new_Sorter100|9736_  | \new_Sorter100|9737_ ;
  assign \new_Sorter100|9838_  = \new_Sorter100|9738_  & \new_Sorter100|9739_ ;
  assign \new_Sorter100|9839_  = \new_Sorter100|9738_  | \new_Sorter100|9739_ ;
  assign \new_Sorter100|9840_  = \new_Sorter100|9740_  & \new_Sorter100|9741_ ;
  assign \new_Sorter100|9841_  = \new_Sorter100|9740_  | \new_Sorter100|9741_ ;
  assign \new_Sorter100|9842_  = \new_Sorter100|9742_  & \new_Sorter100|9743_ ;
  assign \new_Sorter100|9843_  = \new_Sorter100|9742_  | \new_Sorter100|9743_ ;
  assign \new_Sorter100|9844_  = \new_Sorter100|9744_  & \new_Sorter100|9745_ ;
  assign \new_Sorter100|9845_  = \new_Sorter100|9744_  | \new_Sorter100|9745_ ;
  assign \new_Sorter100|9846_  = \new_Sorter100|9746_  & \new_Sorter100|9747_ ;
  assign \new_Sorter100|9847_  = \new_Sorter100|9746_  | \new_Sorter100|9747_ ;
  assign \new_Sorter100|9848_  = \new_Sorter100|9748_  & \new_Sorter100|9749_ ;
  assign \new_Sorter100|9849_  = \new_Sorter100|9748_  | \new_Sorter100|9749_ ;
  assign \new_Sorter100|9850_  = \new_Sorter100|9750_  & \new_Sorter100|9751_ ;
  assign \new_Sorter100|9851_  = \new_Sorter100|9750_  | \new_Sorter100|9751_ ;
  assign \new_Sorter100|9852_  = \new_Sorter100|9752_  & \new_Sorter100|9753_ ;
  assign \new_Sorter100|9853_  = \new_Sorter100|9752_  | \new_Sorter100|9753_ ;
  assign \new_Sorter100|9854_  = \new_Sorter100|9754_  & \new_Sorter100|9755_ ;
  assign \new_Sorter100|9855_  = \new_Sorter100|9754_  | \new_Sorter100|9755_ ;
  assign \new_Sorter100|9856_  = \new_Sorter100|9756_  & \new_Sorter100|9757_ ;
  assign \new_Sorter100|9857_  = \new_Sorter100|9756_  | \new_Sorter100|9757_ ;
  assign \new_Sorter100|9858_  = \new_Sorter100|9758_  & \new_Sorter100|9759_ ;
  assign \new_Sorter100|9859_  = \new_Sorter100|9758_  | \new_Sorter100|9759_ ;
  assign \new_Sorter100|9860_  = \new_Sorter100|9760_  & \new_Sorter100|9761_ ;
  assign \new_Sorter100|9861_  = \new_Sorter100|9760_  | \new_Sorter100|9761_ ;
  assign \new_Sorter100|9862_  = \new_Sorter100|9762_  & \new_Sorter100|9763_ ;
  assign \new_Sorter100|9863_  = \new_Sorter100|9762_  | \new_Sorter100|9763_ ;
  assign \new_Sorter100|9864_  = \new_Sorter100|9764_  & \new_Sorter100|9765_ ;
  assign \new_Sorter100|9865_  = \new_Sorter100|9764_  | \new_Sorter100|9765_ ;
  assign \new_Sorter100|9866_  = \new_Sorter100|9766_  & \new_Sorter100|9767_ ;
  assign \new_Sorter100|9867_  = \new_Sorter100|9766_  | \new_Sorter100|9767_ ;
  assign \new_Sorter100|9868_  = \new_Sorter100|9768_  & \new_Sorter100|9769_ ;
  assign \new_Sorter100|9869_  = \new_Sorter100|9768_  | \new_Sorter100|9769_ ;
  assign \new_Sorter100|9870_  = \new_Sorter100|9770_  & \new_Sorter100|9771_ ;
  assign \new_Sorter100|9871_  = \new_Sorter100|9770_  | \new_Sorter100|9771_ ;
  assign \new_Sorter100|9872_  = \new_Sorter100|9772_  & \new_Sorter100|9773_ ;
  assign \new_Sorter100|9873_  = \new_Sorter100|9772_  | \new_Sorter100|9773_ ;
  assign \new_Sorter100|9874_  = \new_Sorter100|9774_  & \new_Sorter100|9775_ ;
  assign \new_Sorter100|9875_  = \new_Sorter100|9774_  | \new_Sorter100|9775_ ;
  assign \new_Sorter100|9876_  = \new_Sorter100|9776_  & \new_Sorter100|9777_ ;
  assign \new_Sorter100|9877_  = \new_Sorter100|9776_  | \new_Sorter100|9777_ ;
  assign \new_Sorter100|9878_  = \new_Sorter100|9778_  & \new_Sorter100|9779_ ;
  assign \new_Sorter100|9879_  = \new_Sorter100|9778_  | \new_Sorter100|9779_ ;
  assign \new_Sorter100|9880_  = \new_Sorter100|9780_  & \new_Sorter100|9781_ ;
  assign \new_Sorter100|9881_  = \new_Sorter100|9780_  | \new_Sorter100|9781_ ;
  assign \new_Sorter100|9882_  = \new_Sorter100|9782_  & \new_Sorter100|9783_ ;
  assign \new_Sorter100|9883_  = \new_Sorter100|9782_  | \new_Sorter100|9783_ ;
  assign \new_Sorter100|9884_  = \new_Sorter100|9784_  & \new_Sorter100|9785_ ;
  assign \new_Sorter100|9885_  = \new_Sorter100|9784_  | \new_Sorter100|9785_ ;
  assign \new_Sorter100|9886_  = \new_Sorter100|9786_  & \new_Sorter100|9787_ ;
  assign \new_Sorter100|9887_  = \new_Sorter100|9786_  | \new_Sorter100|9787_ ;
  assign \new_Sorter100|9888_  = \new_Sorter100|9788_  & \new_Sorter100|9789_ ;
  assign \new_Sorter100|9889_  = \new_Sorter100|9788_  | \new_Sorter100|9789_ ;
  assign \new_Sorter100|9890_  = \new_Sorter100|9790_  & \new_Sorter100|9791_ ;
  assign \new_Sorter100|9891_  = \new_Sorter100|9790_  | \new_Sorter100|9791_ ;
  assign \new_Sorter100|9892_  = \new_Sorter100|9792_  & \new_Sorter100|9793_ ;
  assign \new_Sorter100|9893_  = \new_Sorter100|9792_  | \new_Sorter100|9793_ ;
  assign \new_Sorter100|9894_  = \new_Sorter100|9794_  & \new_Sorter100|9795_ ;
  assign \new_Sorter100|9895_  = \new_Sorter100|9794_  | \new_Sorter100|9795_ ;
  assign \new_Sorter100|9896_  = \new_Sorter100|9796_  & \new_Sorter100|9797_ ;
  assign \new_Sorter100|9897_  = \new_Sorter100|9796_  | \new_Sorter100|9797_ ;
  assign \new_Sorter100|9898_  = \new_Sorter100|9798_  & \new_Sorter100|9799_ ;
  assign \new_Sorter100|9899_  = \new_Sorter100|9798_  | \new_Sorter100|9799_ ;
  assign \new_Sorter100|9900_  = \new_Sorter100|9800_ ;
  assign \new_Sorter100|9999_  = \new_Sorter100|9899_ ;
  assign \new_Sorter100|9901_  = \new_Sorter100|9801_  & \new_Sorter100|9802_ ;
  assign \new_Sorter100|9902_  = \new_Sorter100|9801_  | \new_Sorter100|9802_ ;
  assign \new_Sorter100|9903_  = \new_Sorter100|9803_  & \new_Sorter100|9804_ ;
  assign \new_Sorter100|9904_  = \new_Sorter100|9803_  | \new_Sorter100|9804_ ;
  assign \new_Sorter100|9905_  = \new_Sorter100|9805_  & \new_Sorter100|9806_ ;
  assign \new_Sorter100|9906_  = \new_Sorter100|9805_  | \new_Sorter100|9806_ ;
  assign \new_Sorter100|9907_  = \new_Sorter100|9807_  & \new_Sorter100|9808_ ;
  assign \new_Sorter100|9908_  = \new_Sorter100|9807_  | \new_Sorter100|9808_ ;
  assign \new_Sorter100|9909_  = \new_Sorter100|9809_  & \new_Sorter100|9810_ ;
  assign \new_Sorter100|9910_  = \new_Sorter100|9809_  | \new_Sorter100|9810_ ;
  assign \new_Sorter100|9911_  = \new_Sorter100|9811_  & \new_Sorter100|9812_ ;
  assign \new_Sorter100|9912_  = \new_Sorter100|9811_  | \new_Sorter100|9812_ ;
  assign \new_Sorter100|9913_  = \new_Sorter100|9813_  & \new_Sorter100|9814_ ;
  assign \new_Sorter100|9914_  = \new_Sorter100|9813_  | \new_Sorter100|9814_ ;
  assign \new_Sorter100|9915_  = \new_Sorter100|9815_  & \new_Sorter100|9816_ ;
  assign \new_Sorter100|9916_  = \new_Sorter100|9815_  | \new_Sorter100|9816_ ;
  assign \new_Sorter100|9917_  = \new_Sorter100|9817_  & \new_Sorter100|9818_ ;
  assign \new_Sorter100|9918_  = \new_Sorter100|9817_  | \new_Sorter100|9818_ ;
  assign \new_Sorter100|9919_  = \new_Sorter100|9819_  & \new_Sorter100|9820_ ;
  assign \new_Sorter100|9920_  = \new_Sorter100|9819_  | \new_Sorter100|9820_ ;
  assign \new_Sorter100|9921_  = \new_Sorter100|9821_  & \new_Sorter100|9822_ ;
  assign \new_Sorter100|9922_  = \new_Sorter100|9821_  | \new_Sorter100|9822_ ;
  assign \new_Sorter100|9923_  = \new_Sorter100|9823_  & \new_Sorter100|9824_ ;
  assign \new_Sorter100|9924_  = \new_Sorter100|9823_  | \new_Sorter100|9824_ ;
  assign \new_Sorter100|9925_  = \new_Sorter100|9825_  & \new_Sorter100|9826_ ;
  assign \new_Sorter100|9926_  = \new_Sorter100|9825_  | \new_Sorter100|9826_ ;
  assign \new_Sorter100|9927_  = \new_Sorter100|9827_  & \new_Sorter100|9828_ ;
  assign \new_Sorter100|9928_  = \new_Sorter100|9827_  | \new_Sorter100|9828_ ;
  assign \new_Sorter100|9929_  = \new_Sorter100|9829_  & \new_Sorter100|9830_ ;
  assign \new_Sorter100|9930_  = \new_Sorter100|9829_  | \new_Sorter100|9830_ ;
  assign \new_Sorter100|9931_  = \new_Sorter100|9831_  & \new_Sorter100|9832_ ;
  assign \new_Sorter100|9932_  = \new_Sorter100|9831_  | \new_Sorter100|9832_ ;
  assign \new_Sorter100|9933_  = \new_Sorter100|9833_  & \new_Sorter100|9834_ ;
  assign \new_Sorter100|9934_  = \new_Sorter100|9833_  | \new_Sorter100|9834_ ;
  assign \new_Sorter100|9935_  = \new_Sorter100|9835_  & \new_Sorter100|9836_ ;
  assign \new_Sorter100|9936_  = \new_Sorter100|9835_  | \new_Sorter100|9836_ ;
  assign \new_Sorter100|9937_  = \new_Sorter100|9837_  & \new_Sorter100|9838_ ;
  assign \new_Sorter100|9938_  = \new_Sorter100|9837_  | \new_Sorter100|9838_ ;
  assign \new_Sorter100|9939_  = \new_Sorter100|9839_  & \new_Sorter100|9840_ ;
  assign \new_Sorter100|9940_  = \new_Sorter100|9839_  | \new_Sorter100|9840_ ;
  assign \new_Sorter100|9941_  = \new_Sorter100|9841_  & \new_Sorter100|9842_ ;
  assign \new_Sorter100|9942_  = \new_Sorter100|9841_  | \new_Sorter100|9842_ ;
  assign \new_Sorter100|9943_  = \new_Sorter100|9843_  & \new_Sorter100|9844_ ;
  assign \new_Sorter100|9944_  = \new_Sorter100|9843_  | \new_Sorter100|9844_ ;
  assign \new_Sorter100|9945_  = \new_Sorter100|9845_  & \new_Sorter100|9846_ ;
  assign \new_Sorter100|9946_  = \new_Sorter100|9845_  | \new_Sorter100|9846_ ;
  assign \new_Sorter100|9947_  = \new_Sorter100|9847_  & \new_Sorter100|9848_ ;
  assign \new_Sorter100|9948_  = \new_Sorter100|9847_  | \new_Sorter100|9848_ ;
  assign \new_Sorter100|9949_  = \new_Sorter100|9849_  & \new_Sorter100|9850_ ;
  assign \new_Sorter100|9950_  = \new_Sorter100|9849_  | \new_Sorter100|9850_ ;
  assign \new_Sorter100|9951_  = \new_Sorter100|9851_  & \new_Sorter100|9852_ ;
  assign \new_Sorter100|9952_  = \new_Sorter100|9851_  | \new_Sorter100|9852_ ;
  assign \new_Sorter100|9953_  = \new_Sorter100|9853_  & \new_Sorter100|9854_ ;
  assign \new_Sorter100|9954_  = \new_Sorter100|9853_  | \new_Sorter100|9854_ ;
  assign \new_Sorter100|9955_  = \new_Sorter100|9855_  & \new_Sorter100|9856_ ;
  assign \new_Sorter100|9956_  = \new_Sorter100|9855_  | \new_Sorter100|9856_ ;
  assign \new_Sorter100|9957_  = \new_Sorter100|9857_  & \new_Sorter100|9858_ ;
  assign \new_Sorter100|9958_  = \new_Sorter100|9857_  | \new_Sorter100|9858_ ;
  assign \new_Sorter100|9959_  = \new_Sorter100|9859_  & \new_Sorter100|9860_ ;
  assign \new_Sorter100|9960_  = \new_Sorter100|9859_  | \new_Sorter100|9860_ ;
  assign \new_Sorter100|9961_  = \new_Sorter100|9861_  & \new_Sorter100|9862_ ;
  assign \new_Sorter100|9962_  = \new_Sorter100|9861_  | \new_Sorter100|9862_ ;
  assign \new_Sorter100|9963_  = \new_Sorter100|9863_  & \new_Sorter100|9864_ ;
  assign \new_Sorter100|9964_  = \new_Sorter100|9863_  | \new_Sorter100|9864_ ;
  assign \new_Sorter100|9965_  = \new_Sorter100|9865_  & \new_Sorter100|9866_ ;
  assign \new_Sorter100|9966_  = \new_Sorter100|9865_  | \new_Sorter100|9866_ ;
  assign \new_Sorter100|9967_  = \new_Sorter100|9867_  & \new_Sorter100|9868_ ;
  assign \new_Sorter100|9968_  = \new_Sorter100|9867_  | \new_Sorter100|9868_ ;
  assign \new_Sorter100|9969_  = \new_Sorter100|9869_  & \new_Sorter100|9870_ ;
  assign \new_Sorter100|9970_  = \new_Sorter100|9869_  | \new_Sorter100|9870_ ;
  assign \new_Sorter100|9971_  = \new_Sorter100|9871_  & \new_Sorter100|9872_ ;
  assign \new_Sorter100|9972_  = \new_Sorter100|9871_  | \new_Sorter100|9872_ ;
  assign \new_Sorter100|9973_  = \new_Sorter100|9873_  & \new_Sorter100|9874_ ;
  assign \new_Sorter100|9974_  = \new_Sorter100|9873_  | \new_Sorter100|9874_ ;
  assign \new_Sorter100|9975_  = \new_Sorter100|9875_  & \new_Sorter100|9876_ ;
  assign \new_Sorter100|9976_  = \new_Sorter100|9875_  | \new_Sorter100|9876_ ;
  assign \new_Sorter100|9977_  = \new_Sorter100|9877_  & \new_Sorter100|9878_ ;
  assign \new_Sorter100|9978_  = \new_Sorter100|9877_  | \new_Sorter100|9878_ ;
  assign \new_Sorter100|9979_  = \new_Sorter100|9879_  & \new_Sorter100|9880_ ;
  assign \new_Sorter100|9980_  = \new_Sorter100|9879_  | \new_Sorter100|9880_ ;
  assign \new_Sorter100|9981_  = \new_Sorter100|9881_  & \new_Sorter100|9882_ ;
  assign \new_Sorter100|9982_  = \new_Sorter100|9881_  | \new_Sorter100|9882_ ;
  assign \new_Sorter100|9983_  = \new_Sorter100|9883_  & \new_Sorter100|9884_ ;
  assign \new_Sorter100|9984_  = \new_Sorter100|9883_  | \new_Sorter100|9884_ ;
  assign \new_Sorter100|9985_  = \new_Sorter100|9885_  & \new_Sorter100|9886_ ;
  assign \new_Sorter100|9986_  = \new_Sorter100|9885_  | \new_Sorter100|9886_ ;
  assign \new_Sorter100|9987_  = \new_Sorter100|9887_  & \new_Sorter100|9888_ ;
  assign \new_Sorter100|9988_  = \new_Sorter100|9887_  | \new_Sorter100|9888_ ;
  assign \new_Sorter100|9989_  = \new_Sorter100|9889_  & \new_Sorter100|9890_ ;
  assign \new_Sorter100|9990_  = \new_Sorter100|9889_  | \new_Sorter100|9890_ ;
  assign \new_Sorter100|9991_  = \new_Sorter100|9891_  & \new_Sorter100|9892_ ;
  assign \new_Sorter100|9992_  = \new_Sorter100|9891_  | \new_Sorter100|9892_ ;
  assign \new_Sorter100|9993_  = \new_Sorter100|9893_  & \new_Sorter100|9894_ ;
  assign \new_Sorter100|9994_  = \new_Sorter100|9893_  | \new_Sorter100|9894_ ;
  assign \new_Sorter100|9995_  = \new_Sorter100|9895_  & \new_Sorter100|9896_ ;
  assign \new_Sorter100|9996_  = \new_Sorter100|9895_  | \new_Sorter100|9896_ ;
  assign \new_Sorter100|9997_  = \new_Sorter100|9897_  & \new_Sorter100|9898_ ;
  assign \new_Sorter100|9998_  = \new_Sorter100|9897_  | \new_Sorter100|9898_ ;
  assign \new_Sorter100|10000_  = \new_Sorter100|9900_  & \new_Sorter100|9901_ ;
  assign \new_Sorter100|10001_  = \new_Sorter100|9900_  | \new_Sorter100|9901_ ;
  assign \new_Sorter100|10002_  = \new_Sorter100|9902_  & \new_Sorter100|9903_ ;
  assign \new_Sorter100|10003_  = \new_Sorter100|9902_  | \new_Sorter100|9903_ ;
  assign \new_Sorter100|10004_  = \new_Sorter100|9904_  & \new_Sorter100|9905_ ;
  assign \new_Sorter100|10005_  = \new_Sorter100|9904_  | \new_Sorter100|9905_ ;
  assign \new_Sorter100|10006_  = \new_Sorter100|9906_  & \new_Sorter100|9907_ ;
  assign \new_Sorter100|10007_  = \new_Sorter100|9906_  | \new_Sorter100|9907_ ;
  assign \new_Sorter100|10008_  = \new_Sorter100|9908_  & \new_Sorter100|9909_ ;
  assign \new_Sorter100|10009_  = \new_Sorter100|9908_  | \new_Sorter100|9909_ ;
  assign \new_Sorter100|10010_  = \new_Sorter100|9910_  & \new_Sorter100|9911_ ;
  assign \new_Sorter100|10011_  = \new_Sorter100|9910_  | \new_Sorter100|9911_ ;
  assign \new_Sorter100|10012_  = \new_Sorter100|9912_  & \new_Sorter100|9913_ ;
  assign \new_Sorter100|10013_  = \new_Sorter100|9912_  | \new_Sorter100|9913_ ;
  assign \new_Sorter100|10014_  = \new_Sorter100|9914_  & \new_Sorter100|9915_ ;
  assign \new_Sorter100|10015_  = \new_Sorter100|9914_  | \new_Sorter100|9915_ ;
  assign \new_Sorter100|10016_  = \new_Sorter100|9916_  & \new_Sorter100|9917_ ;
  assign \new_Sorter100|10017_  = \new_Sorter100|9916_  | \new_Sorter100|9917_ ;
  assign \new_Sorter100|10018_  = \new_Sorter100|9918_  & \new_Sorter100|9919_ ;
  assign \new_Sorter100|10019_  = \new_Sorter100|9918_  | \new_Sorter100|9919_ ;
  assign \new_Sorter100|10020_  = \new_Sorter100|9920_  & \new_Sorter100|9921_ ;
  assign \new_Sorter100|10021_  = \new_Sorter100|9920_  | \new_Sorter100|9921_ ;
  assign \new_Sorter100|10022_  = \new_Sorter100|9922_  & \new_Sorter100|9923_ ;
  assign \new_Sorter100|10023_  = \new_Sorter100|9922_  | \new_Sorter100|9923_ ;
  assign \new_Sorter100|10024_  = \new_Sorter100|9924_  & \new_Sorter100|9925_ ;
  assign \new_Sorter100|10025_  = \new_Sorter100|9924_  | \new_Sorter100|9925_ ;
  assign \new_Sorter100|10026_  = \new_Sorter100|9926_  & \new_Sorter100|9927_ ;
  assign \new_Sorter100|10027_  = \new_Sorter100|9926_  | \new_Sorter100|9927_ ;
  assign \new_Sorter100|10028_  = \new_Sorter100|9928_  & \new_Sorter100|9929_ ;
  assign \new_Sorter100|10029_  = \new_Sorter100|9928_  | \new_Sorter100|9929_ ;
  assign \new_Sorter100|10030_  = \new_Sorter100|9930_  & \new_Sorter100|9931_ ;
  assign \new_Sorter100|10031_  = \new_Sorter100|9930_  | \new_Sorter100|9931_ ;
  assign \new_Sorter100|10032_  = \new_Sorter100|9932_  & \new_Sorter100|9933_ ;
  assign \new_Sorter100|10033_  = \new_Sorter100|9932_  | \new_Sorter100|9933_ ;
  assign \new_Sorter100|10034_  = \new_Sorter100|9934_  & \new_Sorter100|9935_ ;
  assign \new_Sorter100|10035_  = \new_Sorter100|9934_  | \new_Sorter100|9935_ ;
  assign \new_Sorter100|10036_  = \new_Sorter100|9936_  & \new_Sorter100|9937_ ;
  assign \new_Sorter100|10037_  = \new_Sorter100|9936_  | \new_Sorter100|9937_ ;
  assign \new_Sorter100|10038_  = \new_Sorter100|9938_  & \new_Sorter100|9939_ ;
  assign \new_Sorter100|10039_  = \new_Sorter100|9938_  | \new_Sorter100|9939_ ;
  assign \new_Sorter100|10040_  = \new_Sorter100|9940_  & \new_Sorter100|9941_ ;
  assign \new_Sorter100|10041_  = \new_Sorter100|9940_  | \new_Sorter100|9941_ ;
  assign \new_Sorter100|10042_  = \new_Sorter100|9942_  & \new_Sorter100|9943_ ;
  assign \new_Sorter100|10043_  = \new_Sorter100|9942_  | \new_Sorter100|9943_ ;
  assign \new_Sorter100|10044_  = \new_Sorter100|9944_  & \new_Sorter100|9945_ ;
  assign \new_Sorter100|10045_  = \new_Sorter100|9944_  | \new_Sorter100|9945_ ;
  assign \new_Sorter100|10046_  = \new_Sorter100|9946_  & \new_Sorter100|9947_ ;
  assign \new_Sorter100|10047_  = \new_Sorter100|9946_  | \new_Sorter100|9947_ ;
  assign \new_Sorter100|10048_  = \new_Sorter100|9948_  & \new_Sorter100|9949_ ;
  assign \new_Sorter100|10049_  = \new_Sorter100|9948_  | \new_Sorter100|9949_ ;
  assign \new_Sorter100|10050_  = \new_Sorter100|9950_  & \new_Sorter100|9951_ ;
  assign \new_Sorter100|10051_  = \new_Sorter100|9950_  | \new_Sorter100|9951_ ;
  assign \new_Sorter100|10052_  = \new_Sorter100|9952_  & \new_Sorter100|9953_ ;
  assign \new_Sorter100|10053_  = \new_Sorter100|9952_  | \new_Sorter100|9953_ ;
  assign \new_Sorter100|10054_  = \new_Sorter100|9954_  & \new_Sorter100|9955_ ;
  assign \new_Sorter100|10055_  = \new_Sorter100|9954_  | \new_Sorter100|9955_ ;
  assign \new_Sorter100|10056_  = \new_Sorter100|9956_  & \new_Sorter100|9957_ ;
  assign \new_Sorter100|10057_  = \new_Sorter100|9956_  | \new_Sorter100|9957_ ;
  assign \new_Sorter100|10058_  = \new_Sorter100|9958_  & \new_Sorter100|9959_ ;
  assign \new_Sorter100|10059_  = \new_Sorter100|9958_  | \new_Sorter100|9959_ ;
  assign \new_Sorter100|10060_  = \new_Sorter100|9960_  & \new_Sorter100|9961_ ;
  assign \new_Sorter100|10061_  = \new_Sorter100|9960_  | \new_Sorter100|9961_ ;
  assign \new_Sorter100|10062_  = \new_Sorter100|9962_  & \new_Sorter100|9963_ ;
  assign \new_Sorter100|10063_  = \new_Sorter100|9962_  | \new_Sorter100|9963_ ;
  assign \new_Sorter100|10064_  = \new_Sorter100|9964_  & \new_Sorter100|9965_ ;
  assign \new_Sorter100|10065_  = \new_Sorter100|9964_  | \new_Sorter100|9965_ ;
  assign \new_Sorter100|10066_  = \new_Sorter100|9966_  & \new_Sorter100|9967_ ;
  assign \new_Sorter100|10067_  = \new_Sorter100|9966_  | \new_Sorter100|9967_ ;
  assign \new_Sorter100|10068_  = \new_Sorter100|9968_  & \new_Sorter100|9969_ ;
  assign \new_Sorter100|10069_  = \new_Sorter100|9968_  | \new_Sorter100|9969_ ;
  assign \new_Sorter100|10070_  = \new_Sorter100|9970_  & \new_Sorter100|9971_ ;
  assign \new_Sorter100|10071_  = \new_Sorter100|9970_  | \new_Sorter100|9971_ ;
  assign \new_Sorter100|10072_  = \new_Sorter100|9972_  & \new_Sorter100|9973_ ;
  assign \new_Sorter100|10073_  = \new_Sorter100|9972_  | \new_Sorter100|9973_ ;
  assign \new_Sorter100|10074_  = \new_Sorter100|9974_  & \new_Sorter100|9975_ ;
  assign \new_Sorter100|10075_  = \new_Sorter100|9974_  | \new_Sorter100|9975_ ;
  assign \new_Sorter100|10076_  = \new_Sorter100|9976_  & \new_Sorter100|9977_ ;
  assign \new_Sorter100|10077_  = \new_Sorter100|9976_  | \new_Sorter100|9977_ ;
  assign \new_Sorter100|10078_  = \new_Sorter100|9978_  & \new_Sorter100|9979_ ;
  assign \new_Sorter100|10079_  = \new_Sorter100|9978_  | \new_Sorter100|9979_ ;
  assign \new_Sorter100|10080_  = \new_Sorter100|9980_  & \new_Sorter100|9981_ ;
  assign \new_Sorter100|10081_  = \new_Sorter100|9980_  | \new_Sorter100|9981_ ;
  assign \new_Sorter100|10082_  = \new_Sorter100|9982_  & \new_Sorter100|9983_ ;
  assign \new_Sorter100|10083_  = \new_Sorter100|9982_  | \new_Sorter100|9983_ ;
  assign \new_Sorter100|10084_  = \new_Sorter100|9984_  & \new_Sorter100|9985_ ;
  assign \new_Sorter100|10085_  = \new_Sorter100|9984_  | \new_Sorter100|9985_ ;
  assign \new_Sorter100|10086_  = \new_Sorter100|9986_  & \new_Sorter100|9987_ ;
  assign \new_Sorter100|10087_  = \new_Sorter100|9986_  | \new_Sorter100|9987_ ;
  assign \new_Sorter100|10088_  = \new_Sorter100|9988_  & \new_Sorter100|9989_ ;
  assign \new_Sorter100|10089_  = \new_Sorter100|9988_  | \new_Sorter100|9989_ ;
  assign \new_Sorter100|10090_  = \new_Sorter100|9990_  & \new_Sorter100|9991_ ;
  assign \new_Sorter100|10091_  = \new_Sorter100|9990_  | \new_Sorter100|9991_ ;
  assign \new_Sorter100|10092_  = \new_Sorter100|9992_  & \new_Sorter100|9993_ ;
  assign \new_Sorter100|10093_  = \new_Sorter100|9992_  | \new_Sorter100|9993_ ;
  assign \new_Sorter100|10094_  = \new_Sorter100|9994_  & \new_Sorter100|9995_ ;
  assign \new_Sorter100|10095_  = \new_Sorter100|9994_  | \new_Sorter100|9995_ ;
  assign \new_Sorter100|10096_  = \new_Sorter100|9996_  & \new_Sorter100|9997_ ;
  assign \new_Sorter100|10097_  = \new_Sorter100|9996_  | \new_Sorter100|9997_ ;
  assign \new_Sorter100|10098_  = \new_Sorter100|9998_  & \new_Sorter100|9999_ ;
  assign \new_Sorter100|10099_  = \new_Sorter100|9998_  | \new_Sorter100|9999_ ;
  assign \new_Sorter100|10100_  = \new_Sorter100|10000_ ;
  assign \new_Sorter100|10199_  = \new_Sorter100|10099_ ;
  assign \new_Sorter100|10101_  = \new_Sorter100|10001_  & \new_Sorter100|10002_ ;
  assign \new_Sorter100|10102_  = \new_Sorter100|10001_  | \new_Sorter100|10002_ ;
  assign \new_Sorter100|10103_  = \new_Sorter100|10003_  & \new_Sorter100|10004_ ;
  assign \new_Sorter100|10104_  = \new_Sorter100|10003_  | \new_Sorter100|10004_ ;
  assign \new_Sorter100|10105_  = \new_Sorter100|10005_  & \new_Sorter100|10006_ ;
  assign \new_Sorter100|10106_  = \new_Sorter100|10005_  | \new_Sorter100|10006_ ;
  assign \new_Sorter100|10107_  = \new_Sorter100|10007_  & \new_Sorter100|10008_ ;
  assign \new_Sorter100|10108_  = \new_Sorter100|10007_  | \new_Sorter100|10008_ ;
  assign \new_Sorter100|10109_  = \new_Sorter100|10009_  & \new_Sorter100|10010_ ;
  assign \new_Sorter100|10110_  = \new_Sorter100|10009_  | \new_Sorter100|10010_ ;
  assign \new_Sorter100|10111_  = \new_Sorter100|10011_  & \new_Sorter100|10012_ ;
  assign \new_Sorter100|10112_  = \new_Sorter100|10011_  | \new_Sorter100|10012_ ;
  assign \new_Sorter100|10113_  = \new_Sorter100|10013_  & \new_Sorter100|10014_ ;
  assign \new_Sorter100|10114_  = \new_Sorter100|10013_  | \new_Sorter100|10014_ ;
  assign \new_Sorter100|10115_  = \new_Sorter100|10015_  & \new_Sorter100|10016_ ;
  assign \new_Sorter100|10116_  = \new_Sorter100|10015_  | \new_Sorter100|10016_ ;
  assign \new_Sorter100|10117_  = \new_Sorter100|10017_  & \new_Sorter100|10018_ ;
  assign \new_Sorter100|10118_  = \new_Sorter100|10017_  | \new_Sorter100|10018_ ;
  assign \new_Sorter100|10119_  = \new_Sorter100|10019_  & \new_Sorter100|10020_ ;
  assign \new_Sorter100|10120_  = \new_Sorter100|10019_  | \new_Sorter100|10020_ ;
  assign \new_Sorter100|10121_  = \new_Sorter100|10021_  & \new_Sorter100|10022_ ;
  assign \new_Sorter100|10122_  = \new_Sorter100|10021_  | \new_Sorter100|10022_ ;
  assign \new_Sorter100|10123_  = \new_Sorter100|10023_  & \new_Sorter100|10024_ ;
  assign \new_Sorter100|10124_  = \new_Sorter100|10023_  | \new_Sorter100|10024_ ;
  assign \new_Sorter100|10125_  = \new_Sorter100|10025_  & \new_Sorter100|10026_ ;
  assign \new_Sorter100|10126_  = \new_Sorter100|10025_  | \new_Sorter100|10026_ ;
  assign \new_Sorter100|10127_  = \new_Sorter100|10027_  & \new_Sorter100|10028_ ;
  assign \new_Sorter100|10128_  = \new_Sorter100|10027_  | \new_Sorter100|10028_ ;
  assign \new_Sorter100|10129_  = \new_Sorter100|10029_  & \new_Sorter100|10030_ ;
  assign \new_Sorter100|10130_  = \new_Sorter100|10029_  | \new_Sorter100|10030_ ;
  assign \new_Sorter100|10131_  = \new_Sorter100|10031_  & \new_Sorter100|10032_ ;
  assign \new_Sorter100|10132_  = \new_Sorter100|10031_  | \new_Sorter100|10032_ ;
  assign \new_Sorter100|10133_  = \new_Sorter100|10033_  & \new_Sorter100|10034_ ;
  assign \new_Sorter100|10134_  = \new_Sorter100|10033_  | \new_Sorter100|10034_ ;
  assign \new_Sorter100|10135_  = \new_Sorter100|10035_  & \new_Sorter100|10036_ ;
  assign \new_Sorter100|10136_  = \new_Sorter100|10035_  | \new_Sorter100|10036_ ;
  assign \new_Sorter100|10137_  = \new_Sorter100|10037_  & \new_Sorter100|10038_ ;
  assign \new_Sorter100|10138_  = \new_Sorter100|10037_  | \new_Sorter100|10038_ ;
  assign \new_Sorter100|10139_  = \new_Sorter100|10039_  & \new_Sorter100|10040_ ;
  assign \new_Sorter100|10140_  = \new_Sorter100|10039_  | \new_Sorter100|10040_ ;
  assign \new_Sorter100|10141_  = \new_Sorter100|10041_  & \new_Sorter100|10042_ ;
  assign \new_Sorter100|10142_  = \new_Sorter100|10041_  | \new_Sorter100|10042_ ;
  assign \new_Sorter100|10143_  = \new_Sorter100|10043_  & \new_Sorter100|10044_ ;
  assign \new_Sorter100|10144_  = \new_Sorter100|10043_  | \new_Sorter100|10044_ ;
  assign \new_Sorter100|10145_  = \new_Sorter100|10045_  & \new_Sorter100|10046_ ;
  assign \new_Sorter100|10146_  = \new_Sorter100|10045_  | \new_Sorter100|10046_ ;
  assign \new_Sorter100|10147_  = \new_Sorter100|10047_  & \new_Sorter100|10048_ ;
  assign \new_Sorter100|10148_  = \new_Sorter100|10047_  | \new_Sorter100|10048_ ;
  assign \new_Sorter100|10149_  = \new_Sorter100|10049_  & \new_Sorter100|10050_ ;
  assign \new_Sorter100|10150_  = \new_Sorter100|10049_  | \new_Sorter100|10050_ ;
  assign \new_Sorter100|10151_  = \new_Sorter100|10051_  & \new_Sorter100|10052_ ;
  assign \new_Sorter100|10152_  = \new_Sorter100|10051_  | \new_Sorter100|10052_ ;
  assign \new_Sorter100|10153_  = \new_Sorter100|10053_  & \new_Sorter100|10054_ ;
  assign \new_Sorter100|10154_  = \new_Sorter100|10053_  | \new_Sorter100|10054_ ;
  assign \new_Sorter100|10155_  = \new_Sorter100|10055_  & \new_Sorter100|10056_ ;
  assign \new_Sorter100|10156_  = \new_Sorter100|10055_  | \new_Sorter100|10056_ ;
  assign \new_Sorter100|10157_  = \new_Sorter100|10057_  & \new_Sorter100|10058_ ;
  assign \new_Sorter100|10158_  = \new_Sorter100|10057_  | \new_Sorter100|10058_ ;
  assign \new_Sorter100|10159_  = \new_Sorter100|10059_  & \new_Sorter100|10060_ ;
  assign \new_Sorter100|10160_  = \new_Sorter100|10059_  | \new_Sorter100|10060_ ;
  assign \new_Sorter100|10161_  = \new_Sorter100|10061_  & \new_Sorter100|10062_ ;
  assign \new_Sorter100|10162_  = \new_Sorter100|10061_  | \new_Sorter100|10062_ ;
  assign \new_Sorter100|10163_  = \new_Sorter100|10063_  & \new_Sorter100|10064_ ;
  assign \new_Sorter100|10164_  = \new_Sorter100|10063_  | \new_Sorter100|10064_ ;
  assign \new_Sorter100|10165_  = \new_Sorter100|10065_  & \new_Sorter100|10066_ ;
  assign \new_Sorter100|10166_  = \new_Sorter100|10065_  | \new_Sorter100|10066_ ;
  assign \new_Sorter100|10167_  = \new_Sorter100|10067_  & \new_Sorter100|10068_ ;
  assign \new_Sorter100|10168_  = \new_Sorter100|10067_  | \new_Sorter100|10068_ ;
  assign \new_Sorter100|10169_  = \new_Sorter100|10069_  & \new_Sorter100|10070_ ;
  assign \new_Sorter100|10170_  = \new_Sorter100|10069_  | \new_Sorter100|10070_ ;
  assign \new_Sorter100|10171_  = \new_Sorter100|10071_  & \new_Sorter100|10072_ ;
  assign \new_Sorter100|10172_  = \new_Sorter100|10071_  | \new_Sorter100|10072_ ;
  assign \new_Sorter100|10173_  = \new_Sorter100|10073_  & \new_Sorter100|10074_ ;
  assign \new_Sorter100|10174_  = \new_Sorter100|10073_  | \new_Sorter100|10074_ ;
  assign \new_Sorter100|10175_  = \new_Sorter100|10075_  & \new_Sorter100|10076_ ;
  assign \new_Sorter100|10176_  = \new_Sorter100|10075_  | \new_Sorter100|10076_ ;
  assign \new_Sorter100|10177_  = \new_Sorter100|10077_  & \new_Sorter100|10078_ ;
  assign \new_Sorter100|10178_  = \new_Sorter100|10077_  | \new_Sorter100|10078_ ;
  assign \new_Sorter100|10179_  = \new_Sorter100|10079_  & \new_Sorter100|10080_ ;
  assign \new_Sorter100|10180_  = \new_Sorter100|10079_  | \new_Sorter100|10080_ ;
  assign \new_Sorter100|10181_  = \new_Sorter100|10081_  & \new_Sorter100|10082_ ;
  assign \new_Sorter100|10182_  = \new_Sorter100|10081_  | \new_Sorter100|10082_ ;
  assign \new_Sorter100|10183_  = \new_Sorter100|10083_  & \new_Sorter100|10084_ ;
  assign \new_Sorter100|10184_  = \new_Sorter100|10083_  | \new_Sorter100|10084_ ;
  assign \new_Sorter100|10185_  = \new_Sorter100|10085_  & \new_Sorter100|10086_ ;
  assign \new_Sorter100|10186_  = \new_Sorter100|10085_  | \new_Sorter100|10086_ ;
  assign \new_Sorter100|10187_  = \new_Sorter100|10087_  & \new_Sorter100|10088_ ;
  assign \new_Sorter100|10188_  = \new_Sorter100|10087_  | \new_Sorter100|10088_ ;
  assign \new_Sorter100|10189_  = \new_Sorter100|10089_  & \new_Sorter100|10090_ ;
  assign \new_Sorter100|10190_  = \new_Sorter100|10089_  | \new_Sorter100|10090_ ;
  assign \new_Sorter100|10191_  = \new_Sorter100|10091_  & \new_Sorter100|10092_ ;
  assign \new_Sorter100|10192_  = \new_Sorter100|10091_  | \new_Sorter100|10092_ ;
  assign \new_Sorter100|10193_  = \new_Sorter100|10093_  & \new_Sorter100|10094_ ;
  assign \new_Sorter100|10194_  = \new_Sorter100|10093_  | \new_Sorter100|10094_ ;
  assign \new_Sorter100|10195_  = \new_Sorter100|10095_  & \new_Sorter100|10096_ ;
  assign \new_Sorter100|10196_  = \new_Sorter100|10095_  | \new_Sorter100|10096_ ;
  assign \new_Sorter100|10197_  = \new_Sorter100|10097_  & \new_Sorter100|10098_ ;
  assign \new_Sorter100|10198_  = \new_Sorter100|10097_  | \new_Sorter100|10098_ ;
  assign \new_Sorter100|10200_  = \new_Sorter100|10100_  & \new_Sorter100|10101_ ;
  assign \new_Sorter100|10201_  = \new_Sorter100|10100_  | \new_Sorter100|10101_ ;
  assign \new_Sorter100|10202_  = \new_Sorter100|10102_  & \new_Sorter100|10103_ ;
  assign \new_Sorter100|10203_  = \new_Sorter100|10102_  | \new_Sorter100|10103_ ;
  assign \new_Sorter100|10204_  = \new_Sorter100|10104_  & \new_Sorter100|10105_ ;
  assign \new_Sorter100|10205_  = \new_Sorter100|10104_  | \new_Sorter100|10105_ ;
  assign \new_Sorter100|10206_  = \new_Sorter100|10106_  & \new_Sorter100|10107_ ;
  assign \new_Sorter100|10207_  = \new_Sorter100|10106_  | \new_Sorter100|10107_ ;
  assign \new_Sorter100|10208_  = \new_Sorter100|10108_  & \new_Sorter100|10109_ ;
  assign \new_Sorter100|10209_  = \new_Sorter100|10108_  | \new_Sorter100|10109_ ;
  assign \new_Sorter100|10210_  = \new_Sorter100|10110_  & \new_Sorter100|10111_ ;
  assign \new_Sorter100|10211_  = \new_Sorter100|10110_  | \new_Sorter100|10111_ ;
  assign \new_Sorter100|10212_  = \new_Sorter100|10112_  & \new_Sorter100|10113_ ;
  assign \new_Sorter100|10213_  = \new_Sorter100|10112_  | \new_Sorter100|10113_ ;
  assign \new_Sorter100|10214_  = \new_Sorter100|10114_  & \new_Sorter100|10115_ ;
  assign \new_Sorter100|10215_  = \new_Sorter100|10114_  | \new_Sorter100|10115_ ;
  assign \new_Sorter100|10216_  = \new_Sorter100|10116_  & \new_Sorter100|10117_ ;
  assign \new_Sorter100|10217_  = \new_Sorter100|10116_  | \new_Sorter100|10117_ ;
  assign \new_Sorter100|10218_  = \new_Sorter100|10118_  & \new_Sorter100|10119_ ;
  assign \new_Sorter100|10219_  = \new_Sorter100|10118_  | \new_Sorter100|10119_ ;
  assign \new_Sorter100|10220_  = \new_Sorter100|10120_  & \new_Sorter100|10121_ ;
  assign \new_Sorter100|10221_  = \new_Sorter100|10120_  | \new_Sorter100|10121_ ;
  assign \new_Sorter100|10222_  = \new_Sorter100|10122_  & \new_Sorter100|10123_ ;
  assign \new_Sorter100|10223_  = \new_Sorter100|10122_  | \new_Sorter100|10123_ ;
  assign \new_Sorter100|10224_  = \new_Sorter100|10124_  & \new_Sorter100|10125_ ;
  assign \new_Sorter100|10225_  = \new_Sorter100|10124_  | \new_Sorter100|10125_ ;
  assign \new_Sorter100|10226_  = \new_Sorter100|10126_  & \new_Sorter100|10127_ ;
  assign \new_Sorter100|10227_  = \new_Sorter100|10126_  | \new_Sorter100|10127_ ;
  assign \new_Sorter100|10228_  = \new_Sorter100|10128_  & \new_Sorter100|10129_ ;
  assign \new_Sorter100|10229_  = \new_Sorter100|10128_  | \new_Sorter100|10129_ ;
  assign \new_Sorter100|10230_  = \new_Sorter100|10130_  & \new_Sorter100|10131_ ;
  assign \new_Sorter100|10231_  = \new_Sorter100|10130_  | \new_Sorter100|10131_ ;
  assign \new_Sorter100|10232_  = \new_Sorter100|10132_  & \new_Sorter100|10133_ ;
  assign \new_Sorter100|10233_  = \new_Sorter100|10132_  | \new_Sorter100|10133_ ;
  assign \new_Sorter100|10234_  = \new_Sorter100|10134_  & \new_Sorter100|10135_ ;
  assign \new_Sorter100|10235_  = \new_Sorter100|10134_  | \new_Sorter100|10135_ ;
  assign \new_Sorter100|10236_  = \new_Sorter100|10136_  & \new_Sorter100|10137_ ;
  assign \new_Sorter100|10237_  = \new_Sorter100|10136_  | \new_Sorter100|10137_ ;
  assign \new_Sorter100|10238_  = \new_Sorter100|10138_  & \new_Sorter100|10139_ ;
  assign \new_Sorter100|10239_  = \new_Sorter100|10138_  | \new_Sorter100|10139_ ;
  assign \new_Sorter100|10240_  = \new_Sorter100|10140_  & \new_Sorter100|10141_ ;
  assign \new_Sorter100|10241_  = \new_Sorter100|10140_  | \new_Sorter100|10141_ ;
  assign \new_Sorter100|10242_  = \new_Sorter100|10142_  & \new_Sorter100|10143_ ;
  assign \new_Sorter100|10243_  = \new_Sorter100|10142_  | \new_Sorter100|10143_ ;
  assign \new_Sorter100|10244_  = \new_Sorter100|10144_  & \new_Sorter100|10145_ ;
  assign \new_Sorter100|10245_  = \new_Sorter100|10144_  | \new_Sorter100|10145_ ;
  assign \new_Sorter100|10246_  = \new_Sorter100|10146_  & \new_Sorter100|10147_ ;
  assign \new_Sorter100|10247_  = \new_Sorter100|10146_  | \new_Sorter100|10147_ ;
  assign \new_Sorter100|10248_  = \new_Sorter100|10148_  & \new_Sorter100|10149_ ;
  assign \new_Sorter100|10249_  = \new_Sorter100|10148_  | \new_Sorter100|10149_ ;
  assign \new_Sorter100|10250_  = \new_Sorter100|10150_  & \new_Sorter100|10151_ ;
  assign \new_Sorter100|10251_  = \new_Sorter100|10150_  | \new_Sorter100|10151_ ;
  assign \new_Sorter100|10252_  = \new_Sorter100|10152_  & \new_Sorter100|10153_ ;
  assign \new_Sorter100|10253_  = \new_Sorter100|10152_  | \new_Sorter100|10153_ ;
  assign \new_Sorter100|10254_  = \new_Sorter100|10154_  & \new_Sorter100|10155_ ;
  assign \new_Sorter100|10255_  = \new_Sorter100|10154_  | \new_Sorter100|10155_ ;
  assign \new_Sorter100|10256_  = \new_Sorter100|10156_  & \new_Sorter100|10157_ ;
  assign \new_Sorter100|10257_  = \new_Sorter100|10156_  | \new_Sorter100|10157_ ;
  assign \new_Sorter100|10258_  = \new_Sorter100|10158_  & \new_Sorter100|10159_ ;
  assign \new_Sorter100|10259_  = \new_Sorter100|10158_  | \new_Sorter100|10159_ ;
  assign \new_Sorter100|10260_  = \new_Sorter100|10160_  & \new_Sorter100|10161_ ;
  assign \new_Sorter100|10261_  = \new_Sorter100|10160_  | \new_Sorter100|10161_ ;
  assign \new_Sorter100|10262_  = \new_Sorter100|10162_  & \new_Sorter100|10163_ ;
  assign \new_Sorter100|10263_  = \new_Sorter100|10162_  | \new_Sorter100|10163_ ;
  assign \new_Sorter100|10264_  = \new_Sorter100|10164_  & \new_Sorter100|10165_ ;
  assign \new_Sorter100|10265_  = \new_Sorter100|10164_  | \new_Sorter100|10165_ ;
  assign \new_Sorter100|10266_  = \new_Sorter100|10166_  & \new_Sorter100|10167_ ;
  assign \new_Sorter100|10267_  = \new_Sorter100|10166_  | \new_Sorter100|10167_ ;
  assign \new_Sorter100|10268_  = \new_Sorter100|10168_  & \new_Sorter100|10169_ ;
  assign \new_Sorter100|10269_  = \new_Sorter100|10168_  | \new_Sorter100|10169_ ;
  assign \new_Sorter100|10270_  = \new_Sorter100|10170_  & \new_Sorter100|10171_ ;
  assign \new_Sorter100|10271_  = \new_Sorter100|10170_  | \new_Sorter100|10171_ ;
  assign \new_Sorter100|10272_  = \new_Sorter100|10172_  & \new_Sorter100|10173_ ;
  assign \new_Sorter100|10273_  = \new_Sorter100|10172_  | \new_Sorter100|10173_ ;
  assign \new_Sorter100|10274_  = \new_Sorter100|10174_  & \new_Sorter100|10175_ ;
  assign \new_Sorter100|10275_  = \new_Sorter100|10174_  | \new_Sorter100|10175_ ;
  assign \new_Sorter100|10276_  = \new_Sorter100|10176_  & \new_Sorter100|10177_ ;
  assign \new_Sorter100|10277_  = \new_Sorter100|10176_  | \new_Sorter100|10177_ ;
  assign \new_Sorter100|10278_  = \new_Sorter100|10178_  & \new_Sorter100|10179_ ;
  assign \new_Sorter100|10279_  = \new_Sorter100|10178_  | \new_Sorter100|10179_ ;
  assign \new_Sorter100|10280_  = \new_Sorter100|10180_  & \new_Sorter100|10181_ ;
  assign \new_Sorter100|10281_  = \new_Sorter100|10180_  | \new_Sorter100|10181_ ;
  assign \new_Sorter100|10282_  = \new_Sorter100|10182_  & \new_Sorter100|10183_ ;
  assign \new_Sorter100|10283_  = \new_Sorter100|10182_  | \new_Sorter100|10183_ ;
  assign \new_Sorter100|10284_  = \new_Sorter100|10184_  & \new_Sorter100|10185_ ;
  assign \new_Sorter100|10285_  = \new_Sorter100|10184_  | \new_Sorter100|10185_ ;
  assign \new_Sorter100|10286_  = \new_Sorter100|10186_  & \new_Sorter100|10187_ ;
  assign \new_Sorter100|10287_  = \new_Sorter100|10186_  | \new_Sorter100|10187_ ;
  assign \new_Sorter100|10288_  = \new_Sorter100|10188_  & \new_Sorter100|10189_ ;
  assign \new_Sorter100|10289_  = \new_Sorter100|10188_  | \new_Sorter100|10189_ ;
  assign \new_Sorter100|10290_  = \new_Sorter100|10190_  & \new_Sorter100|10191_ ;
  assign \new_Sorter100|10291_  = \new_Sorter100|10190_  | \new_Sorter100|10191_ ;
  assign \new_Sorter100|10292_  = \new_Sorter100|10192_  & \new_Sorter100|10193_ ;
  assign \new_Sorter100|10293_  = \new_Sorter100|10192_  | \new_Sorter100|10193_ ;
  assign \new_Sorter100|10294_  = \new_Sorter100|10194_  & \new_Sorter100|10195_ ;
  assign \new_Sorter100|10295_  = \new_Sorter100|10194_  | \new_Sorter100|10195_ ;
  assign \new_Sorter100|10296_  = \new_Sorter100|10196_  & \new_Sorter100|10197_ ;
  assign \new_Sorter100|10297_  = \new_Sorter100|10196_  | \new_Sorter100|10197_ ;
  assign \new_Sorter100|10298_  = \new_Sorter100|10198_  & \new_Sorter100|10199_ ;
  assign \new_Sorter100|10299_  = \new_Sorter100|10198_  | \new_Sorter100|10199_ ;
  assign \new_Sorter100|10300_  = \new_Sorter100|10200_ ;
  assign \new_Sorter100|10399_  = \new_Sorter100|10299_ ;
  assign \new_Sorter100|10301_  = \new_Sorter100|10201_  & \new_Sorter100|10202_ ;
  assign \new_Sorter100|10302_  = \new_Sorter100|10201_  | \new_Sorter100|10202_ ;
  assign \new_Sorter100|10303_  = \new_Sorter100|10203_  & \new_Sorter100|10204_ ;
  assign \new_Sorter100|10304_  = \new_Sorter100|10203_  | \new_Sorter100|10204_ ;
  assign \new_Sorter100|10305_  = \new_Sorter100|10205_  & \new_Sorter100|10206_ ;
  assign \new_Sorter100|10306_  = \new_Sorter100|10205_  | \new_Sorter100|10206_ ;
  assign \new_Sorter100|10307_  = \new_Sorter100|10207_  & \new_Sorter100|10208_ ;
  assign \new_Sorter100|10308_  = \new_Sorter100|10207_  | \new_Sorter100|10208_ ;
  assign \new_Sorter100|10309_  = \new_Sorter100|10209_  & \new_Sorter100|10210_ ;
  assign \new_Sorter100|10310_  = \new_Sorter100|10209_  | \new_Sorter100|10210_ ;
  assign \new_Sorter100|10311_  = \new_Sorter100|10211_  & \new_Sorter100|10212_ ;
  assign \new_Sorter100|10312_  = \new_Sorter100|10211_  | \new_Sorter100|10212_ ;
  assign \new_Sorter100|10313_  = \new_Sorter100|10213_  & \new_Sorter100|10214_ ;
  assign \new_Sorter100|10314_  = \new_Sorter100|10213_  | \new_Sorter100|10214_ ;
  assign \new_Sorter100|10315_  = \new_Sorter100|10215_  & \new_Sorter100|10216_ ;
  assign \new_Sorter100|10316_  = \new_Sorter100|10215_  | \new_Sorter100|10216_ ;
  assign \new_Sorter100|10317_  = \new_Sorter100|10217_  & \new_Sorter100|10218_ ;
  assign \new_Sorter100|10318_  = \new_Sorter100|10217_  | \new_Sorter100|10218_ ;
  assign \new_Sorter100|10319_  = \new_Sorter100|10219_  & \new_Sorter100|10220_ ;
  assign \new_Sorter100|10320_  = \new_Sorter100|10219_  | \new_Sorter100|10220_ ;
  assign \new_Sorter100|10321_  = \new_Sorter100|10221_  & \new_Sorter100|10222_ ;
  assign \new_Sorter100|10322_  = \new_Sorter100|10221_  | \new_Sorter100|10222_ ;
  assign \new_Sorter100|10323_  = \new_Sorter100|10223_  & \new_Sorter100|10224_ ;
  assign \new_Sorter100|10324_  = \new_Sorter100|10223_  | \new_Sorter100|10224_ ;
  assign \new_Sorter100|10325_  = \new_Sorter100|10225_  & \new_Sorter100|10226_ ;
  assign \new_Sorter100|10326_  = \new_Sorter100|10225_  | \new_Sorter100|10226_ ;
  assign \new_Sorter100|10327_  = \new_Sorter100|10227_  & \new_Sorter100|10228_ ;
  assign \new_Sorter100|10328_  = \new_Sorter100|10227_  | \new_Sorter100|10228_ ;
  assign \new_Sorter100|10329_  = \new_Sorter100|10229_  & \new_Sorter100|10230_ ;
  assign \new_Sorter100|10330_  = \new_Sorter100|10229_  | \new_Sorter100|10230_ ;
  assign \new_Sorter100|10331_  = \new_Sorter100|10231_  & \new_Sorter100|10232_ ;
  assign \new_Sorter100|10332_  = \new_Sorter100|10231_  | \new_Sorter100|10232_ ;
  assign \new_Sorter100|10333_  = \new_Sorter100|10233_  & \new_Sorter100|10234_ ;
  assign \new_Sorter100|10334_  = \new_Sorter100|10233_  | \new_Sorter100|10234_ ;
  assign \new_Sorter100|10335_  = \new_Sorter100|10235_  & \new_Sorter100|10236_ ;
  assign \new_Sorter100|10336_  = \new_Sorter100|10235_  | \new_Sorter100|10236_ ;
  assign \new_Sorter100|10337_  = \new_Sorter100|10237_  & \new_Sorter100|10238_ ;
  assign \new_Sorter100|10338_  = \new_Sorter100|10237_  | \new_Sorter100|10238_ ;
  assign \new_Sorter100|10339_  = \new_Sorter100|10239_  & \new_Sorter100|10240_ ;
  assign \new_Sorter100|10340_  = \new_Sorter100|10239_  | \new_Sorter100|10240_ ;
  assign \new_Sorter100|10341_  = \new_Sorter100|10241_  & \new_Sorter100|10242_ ;
  assign \new_Sorter100|10342_  = \new_Sorter100|10241_  | \new_Sorter100|10242_ ;
  assign \new_Sorter100|10343_  = \new_Sorter100|10243_  & \new_Sorter100|10244_ ;
  assign \new_Sorter100|10344_  = \new_Sorter100|10243_  | \new_Sorter100|10244_ ;
  assign \new_Sorter100|10345_  = \new_Sorter100|10245_  & \new_Sorter100|10246_ ;
  assign \new_Sorter100|10346_  = \new_Sorter100|10245_  | \new_Sorter100|10246_ ;
  assign \new_Sorter100|10347_  = \new_Sorter100|10247_  & \new_Sorter100|10248_ ;
  assign \new_Sorter100|10348_  = \new_Sorter100|10247_  | \new_Sorter100|10248_ ;
  assign \new_Sorter100|10349_  = \new_Sorter100|10249_  & \new_Sorter100|10250_ ;
  assign \new_Sorter100|10350_  = \new_Sorter100|10249_  | \new_Sorter100|10250_ ;
  assign \new_Sorter100|10351_  = \new_Sorter100|10251_  & \new_Sorter100|10252_ ;
  assign \new_Sorter100|10352_  = \new_Sorter100|10251_  | \new_Sorter100|10252_ ;
  assign \new_Sorter100|10353_  = \new_Sorter100|10253_  & \new_Sorter100|10254_ ;
  assign \new_Sorter100|10354_  = \new_Sorter100|10253_  | \new_Sorter100|10254_ ;
  assign \new_Sorter100|10355_  = \new_Sorter100|10255_  & \new_Sorter100|10256_ ;
  assign \new_Sorter100|10356_  = \new_Sorter100|10255_  | \new_Sorter100|10256_ ;
  assign \new_Sorter100|10357_  = \new_Sorter100|10257_  & \new_Sorter100|10258_ ;
  assign \new_Sorter100|10358_  = \new_Sorter100|10257_  | \new_Sorter100|10258_ ;
  assign \new_Sorter100|10359_  = \new_Sorter100|10259_  & \new_Sorter100|10260_ ;
  assign \new_Sorter100|10360_  = \new_Sorter100|10259_  | \new_Sorter100|10260_ ;
  assign \new_Sorter100|10361_  = \new_Sorter100|10261_  & \new_Sorter100|10262_ ;
  assign \new_Sorter100|10362_  = \new_Sorter100|10261_  | \new_Sorter100|10262_ ;
  assign \new_Sorter100|10363_  = \new_Sorter100|10263_  & \new_Sorter100|10264_ ;
  assign \new_Sorter100|10364_  = \new_Sorter100|10263_  | \new_Sorter100|10264_ ;
  assign \new_Sorter100|10365_  = \new_Sorter100|10265_  & \new_Sorter100|10266_ ;
  assign \new_Sorter100|10366_  = \new_Sorter100|10265_  | \new_Sorter100|10266_ ;
  assign \new_Sorter100|10367_  = \new_Sorter100|10267_  & \new_Sorter100|10268_ ;
  assign \new_Sorter100|10368_  = \new_Sorter100|10267_  | \new_Sorter100|10268_ ;
  assign \new_Sorter100|10369_  = \new_Sorter100|10269_  & \new_Sorter100|10270_ ;
  assign \new_Sorter100|10370_  = \new_Sorter100|10269_  | \new_Sorter100|10270_ ;
  assign \new_Sorter100|10371_  = \new_Sorter100|10271_  & \new_Sorter100|10272_ ;
  assign \new_Sorter100|10372_  = \new_Sorter100|10271_  | \new_Sorter100|10272_ ;
  assign \new_Sorter100|10373_  = \new_Sorter100|10273_  & \new_Sorter100|10274_ ;
  assign \new_Sorter100|10374_  = \new_Sorter100|10273_  | \new_Sorter100|10274_ ;
  assign \new_Sorter100|10375_  = \new_Sorter100|10275_  & \new_Sorter100|10276_ ;
  assign \new_Sorter100|10376_  = \new_Sorter100|10275_  | \new_Sorter100|10276_ ;
  assign \new_Sorter100|10377_  = \new_Sorter100|10277_  & \new_Sorter100|10278_ ;
  assign \new_Sorter100|10378_  = \new_Sorter100|10277_  | \new_Sorter100|10278_ ;
  assign \new_Sorter100|10379_  = \new_Sorter100|10279_  & \new_Sorter100|10280_ ;
  assign \new_Sorter100|10380_  = \new_Sorter100|10279_  | \new_Sorter100|10280_ ;
  assign \new_Sorter100|10381_  = \new_Sorter100|10281_  & \new_Sorter100|10282_ ;
  assign \new_Sorter100|10382_  = \new_Sorter100|10281_  | \new_Sorter100|10282_ ;
  assign \new_Sorter100|10383_  = \new_Sorter100|10283_  & \new_Sorter100|10284_ ;
  assign \new_Sorter100|10384_  = \new_Sorter100|10283_  | \new_Sorter100|10284_ ;
  assign \new_Sorter100|10385_  = \new_Sorter100|10285_  & \new_Sorter100|10286_ ;
  assign \new_Sorter100|10386_  = \new_Sorter100|10285_  | \new_Sorter100|10286_ ;
  assign \new_Sorter100|10387_  = \new_Sorter100|10287_  & \new_Sorter100|10288_ ;
  assign \new_Sorter100|10388_  = \new_Sorter100|10287_  | \new_Sorter100|10288_ ;
  assign \new_Sorter100|10389_  = \new_Sorter100|10289_  & \new_Sorter100|10290_ ;
  assign \new_Sorter100|10390_  = \new_Sorter100|10289_  | \new_Sorter100|10290_ ;
  assign \new_Sorter100|10391_  = \new_Sorter100|10291_  & \new_Sorter100|10292_ ;
  assign \new_Sorter100|10392_  = \new_Sorter100|10291_  | \new_Sorter100|10292_ ;
  assign \new_Sorter100|10393_  = \new_Sorter100|10293_  & \new_Sorter100|10294_ ;
  assign \new_Sorter100|10394_  = \new_Sorter100|10293_  | \new_Sorter100|10294_ ;
  assign \new_Sorter100|10395_  = \new_Sorter100|10295_  & \new_Sorter100|10296_ ;
  assign \new_Sorter100|10396_  = \new_Sorter100|10295_  | \new_Sorter100|10296_ ;
  assign \new_Sorter100|10397_  = \new_Sorter100|10297_  & \new_Sorter100|10298_ ;
  assign \new_Sorter100|10398_  = \new_Sorter100|10297_  | \new_Sorter100|10298_ ;
  assign \new_Sorter100|10400_  = \new_Sorter100|10300_  & \new_Sorter100|10301_ ;
  assign \new_Sorter100|10401_  = \new_Sorter100|10300_  | \new_Sorter100|10301_ ;
  assign \new_Sorter100|10402_  = \new_Sorter100|10302_  & \new_Sorter100|10303_ ;
  assign \new_Sorter100|10403_  = \new_Sorter100|10302_  | \new_Sorter100|10303_ ;
  assign \new_Sorter100|10404_  = \new_Sorter100|10304_  & \new_Sorter100|10305_ ;
  assign \new_Sorter100|10405_  = \new_Sorter100|10304_  | \new_Sorter100|10305_ ;
  assign \new_Sorter100|10406_  = \new_Sorter100|10306_  & \new_Sorter100|10307_ ;
  assign \new_Sorter100|10407_  = \new_Sorter100|10306_  | \new_Sorter100|10307_ ;
  assign \new_Sorter100|10408_  = \new_Sorter100|10308_  & \new_Sorter100|10309_ ;
  assign \new_Sorter100|10409_  = \new_Sorter100|10308_  | \new_Sorter100|10309_ ;
  assign \new_Sorter100|10410_  = \new_Sorter100|10310_  & \new_Sorter100|10311_ ;
  assign \new_Sorter100|10411_  = \new_Sorter100|10310_  | \new_Sorter100|10311_ ;
  assign \new_Sorter100|10412_  = \new_Sorter100|10312_  & \new_Sorter100|10313_ ;
  assign \new_Sorter100|10413_  = \new_Sorter100|10312_  | \new_Sorter100|10313_ ;
  assign \new_Sorter100|10414_  = \new_Sorter100|10314_  & \new_Sorter100|10315_ ;
  assign \new_Sorter100|10415_  = \new_Sorter100|10314_  | \new_Sorter100|10315_ ;
  assign \new_Sorter100|10416_  = \new_Sorter100|10316_  & \new_Sorter100|10317_ ;
  assign \new_Sorter100|10417_  = \new_Sorter100|10316_  | \new_Sorter100|10317_ ;
  assign \new_Sorter100|10418_  = \new_Sorter100|10318_  & \new_Sorter100|10319_ ;
  assign \new_Sorter100|10419_  = \new_Sorter100|10318_  | \new_Sorter100|10319_ ;
  assign \new_Sorter100|10420_  = \new_Sorter100|10320_  & \new_Sorter100|10321_ ;
  assign \new_Sorter100|10421_  = \new_Sorter100|10320_  | \new_Sorter100|10321_ ;
  assign \new_Sorter100|10422_  = \new_Sorter100|10322_  & \new_Sorter100|10323_ ;
  assign \new_Sorter100|10423_  = \new_Sorter100|10322_  | \new_Sorter100|10323_ ;
  assign \new_Sorter100|10424_  = \new_Sorter100|10324_  & \new_Sorter100|10325_ ;
  assign \new_Sorter100|10425_  = \new_Sorter100|10324_  | \new_Sorter100|10325_ ;
  assign \new_Sorter100|10426_  = \new_Sorter100|10326_  & \new_Sorter100|10327_ ;
  assign \new_Sorter100|10427_  = \new_Sorter100|10326_  | \new_Sorter100|10327_ ;
  assign \new_Sorter100|10428_  = \new_Sorter100|10328_  & \new_Sorter100|10329_ ;
  assign \new_Sorter100|10429_  = \new_Sorter100|10328_  | \new_Sorter100|10329_ ;
  assign \new_Sorter100|10430_  = \new_Sorter100|10330_  & \new_Sorter100|10331_ ;
  assign \new_Sorter100|10431_  = \new_Sorter100|10330_  | \new_Sorter100|10331_ ;
  assign \new_Sorter100|10432_  = \new_Sorter100|10332_  & \new_Sorter100|10333_ ;
  assign \new_Sorter100|10433_  = \new_Sorter100|10332_  | \new_Sorter100|10333_ ;
  assign \new_Sorter100|10434_  = \new_Sorter100|10334_  & \new_Sorter100|10335_ ;
  assign \new_Sorter100|10435_  = \new_Sorter100|10334_  | \new_Sorter100|10335_ ;
  assign \new_Sorter100|10436_  = \new_Sorter100|10336_  & \new_Sorter100|10337_ ;
  assign \new_Sorter100|10437_  = \new_Sorter100|10336_  | \new_Sorter100|10337_ ;
  assign \new_Sorter100|10438_  = \new_Sorter100|10338_  & \new_Sorter100|10339_ ;
  assign \new_Sorter100|10439_  = \new_Sorter100|10338_  | \new_Sorter100|10339_ ;
  assign \new_Sorter100|10440_  = \new_Sorter100|10340_  & \new_Sorter100|10341_ ;
  assign \new_Sorter100|10441_  = \new_Sorter100|10340_  | \new_Sorter100|10341_ ;
  assign \new_Sorter100|10442_  = \new_Sorter100|10342_  & \new_Sorter100|10343_ ;
  assign \new_Sorter100|10443_  = \new_Sorter100|10342_  | \new_Sorter100|10343_ ;
  assign \new_Sorter100|10444_  = \new_Sorter100|10344_  & \new_Sorter100|10345_ ;
  assign \new_Sorter100|10445_  = \new_Sorter100|10344_  | \new_Sorter100|10345_ ;
  assign \new_Sorter100|10446_  = \new_Sorter100|10346_  & \new_Sorter100|10347_ ;
  assign \new_Sorter100|10447_  = \new_Sorter100|10346_  | \new_Sorter100|10347_ ;
  assign \new_Sorter100|10448_  = \new_Sorter100|10348_  & \new_Sorter100|10349_ ;
  assign \new_Sorter100|10449_  = \new_Sorter100|10348_  | \new_Sorter100|10349_ ;
  assign \new_Sorter100|10450_  = \new_Sorter100|10350_  & \new_Sorter100|10351_ ;
  assign \new_Sorter100|10451_  = \new_Sorter100|10350_  | \new_Sorter100|10351_ ;
  assign \new_Sorter100|10452_  = \new_Sorter100|10352_  & \new_Sorter100|10353_ ;
  assign \new_Sorter100|10453_  = \new_Sorter100|10352_  | \new_Sorter100|10353_ ;
  assign \new_Sorter100|10454_  = \new_Sorter100|10354_  & \new_Sorter100|10355_ ;
  assign \new_Sorter100|10455_  = \new_Sorter100|10354_  | \new_Sorter100|10355_ ;
  assign \new_Sorter100|10456_  = \new_Sorter100|10356_  & \new_Sorter100|10357_ ;
  assign \new_Sorter100|10457_  = \new_Sorter100|10356_  | \new_Sorter100|10357_ ;
  assign \new_Sorter100|10458_  = \new_Sorter100|10358_  & \new_Sorter100|10359_ ;
  assign \new_Sorter100|10459_  = \new_Sorter100|10358_  | \new_Sorter100|10359_ ;
  assign \new_Sorter100|10460_  = \new_Sorter100|10360_  & \new_Sorter100|10361_ ;
  assign \new_Sorter100|10461_  = \new_Sorter100|10360_  | \new_Sorter100|10361_ ;
  assign \new_Sorter100|10462_  = \new_Sorter100|10362_  & \new_Sorter100|10363_ ;
  assign \new_Sorter100|10463_  = \new_Sorter100|10362_  | \new_Sorter100|10363_ ;
  assign \new_Sorter100|10464_  = \new_Sorter100|10364_  & \new_Sorter100|10365_ ;
  assign \new_Sorter100|10465_  = \new_Sorter100|10364_  | \new_Sorter100|10365_ ;
  assign \new_Sorter100|10466_  = \new_Sorter100|10366_  & \new_Sorter100|10367_ ;
  assign \new_Sorter100|10467_  = \new_Sorter100|10366_  | \new_Sorter100|10367_ ;
  assign \new_Sorter100|10468_  = \new_Sorter100|10368_  & \new_Sorter100|10369_ ;
  assign \new_Sorter100|10469_  = \new_Sorter100|10368_  | \new_Sorter100|10369_ ;
  assign \new_Sorter100|10470_  = \new_Sorter100|10370_  & \new_Sorter100|10371_ ;
  assign \new_Sorter100|10471_  = \new_Sorter100|10370_  | \new_Sorter100|10371_ ;
  assign \new_Sorter100|10472_  = \new_Sorter100|10372_  & \new_Sorter100|10373_ ;
  assign \new_Sorter100|10473_  = \new_Sorter100|10372_  | \new_Sorter100|10373_ ;
  assign \new_Sorter100|10474_  = \new_Sorter100|10374_  & \new_Sorter100|10375_ ;
  assign \new_Sorter100|10475_  = \new_Sorter100|10374_  | \new_Sorter100|10375_ ;
  assign \new_Sorter100|10476_  = \new_Sorter100|10376_  & \new_Sorter100|10377_ ;
  assign \new_Sorter100|10477_  = \new_Sorter100|10376_  | \new_Sorter100|10377_ ;
  assign \new_Sorter100|10478_  = \new_Sorter100|10378_  & \new_Sorter100|10379_ ;
  assign \new_Sorter100|10479_  = \new_Sorter100|10378_  | \new_Sorter100|10379_ ;
  assign \new_Sorter100|10480_  = \new_Sorter100|10380_  & \new_Sorter100|10381_ ;
  assign \new_Sorter100|10481_  = \new_Sorter100|10380_  | \new_Sorter100|10381_ ;
  assign \new_Sorter100|10482_  = \new_Sorter100|10382_  & \new_Sorter100|10383_ ;
  assign \new_Sorter100|10483_  = \new_Sorter100|10382_  | \new_Sorter100|10383_ ;
  assign \new_Sorter100|10484_  = \new_Sorter100|10384_  & \new_Sorter100|10385_ ;
  assign \new_Sorter100|10485_  = \new_Sorter100|10384_  | \new_Sorter100|10385_ ;
  assign \new_Sorter100|10486_  = \new_Sorter100|10386_  & \new_Sorter100|10387_ ;
  assign \new_Sorter100|10487_  = \new_Sorter100|10386_  | \new_Sorter100|10387_ ;
  assign \new_Sorter100|10488_  = \new_Sorter100|10388_  & \new_Sorter100|10389_ ;
  assign \new_Sorter100|10489_  = \new_Sorter100|10388_  | \new_Sorter100|10389_ ;
  assign \new_Sorter100|10490_  = \new_Sorter100|10390_  & \new_Sorter100|10391_ ;
  assign \new_Sorter100|10491_  = \new_Sorter100|10390_  | \new_Sorter100|10391_ ;
  assign \new_Sorter100|10492_  = \new_Sorter100|10392_  & \new_Sorter100|10393_ ;
  assign \new_Sorter100|10493_  = \new_Sorter100|10392_  | \new_Sorter100|10393_ ;
  assign \new_Sorter100|10494_  = \new_Sorter100|10394_  & \new_Sorter100|10395_ ;
  assign \new_Sorter100|10495_  = \new_Sorter100|10394_  | \new_Sorter100|10395_ ;
  assign \new_Sorter100|10496_  = \new_Sorter100|10396_  & \new_Sorter100|10397_ ;
  assign \new_Sorter100|10497_  = \new_Sorter100|10396_  | \new_Sorter100|10397_ ;
  assign \new_Sorter100|10498_  = \new_Sorter100|10398_  & \new_Sorter100|10399_ ;
  assign \new_Sorter100|10499_  = \new_Sorter100|10398_  | \new_Sorter100|10399_ ;
  assign \new_Sorter100|10500_  = \new_Sorter100|10400_ ;
  assign \new_Sorter100|10599_  = \new_Sorter100|10499_ ;
  assign \new_Sorter100|10501_  = \new_Sorter100|10401_  & \new_Sorter100|10402_ ;
  assign \new_Sorter100|10502_  = \new_Sorter100|10401_  | \new_Sorter100|10402_ ;
  assign \new_Sorter100|10503_  = \new_Sorter100|10403_  & \new_Sorter100|10404_ ;
  assign \new_Sorter100|10504_  = \new_Sorter100|10403_  | \new_Sorter100|10404_ ;
  assign \new_Sorter100|10505_  = \new_Sorter100|10405_  & \new_Sorter100|10406_ ;
  assign \new_Sorter100|10506_  = \new_Sorter100|10405_  | \new_Sorter100|10406_ ;
  assign \new_Sorter100|10507_  = \new_Sorter100|10407_  & \new_Sorter100|10408_ ;
  assign \new_Sorter100|10508_  = \new_Sorter100|10407_  | \new_Sorter100|10408_ ;
  assign \new_Sorter100|10509_  = \new_Sorter100|10409_  & \new_Sorter100|10410_ ;
  assign \new_Sorter100|10510_  = \new_Sorter100|10409_  | \new_Sorter100|10410_ ;
  assign \new_Sorter100|10511_  = \new_Sorter100|10411_  & \new_Sorter100|10412_ ;
  assign \new_Sorter100|10512_  = \new_Sorter100|10411_  | \new_Sorter100|10412_ ;
  assign \new_Sorter100|10513_  = \new_Sorter100|10413_  & \new_Sorter100|10414_ ;
  assign \new_Sorter100|10514_  = \new_Sorter100|10413_  | \new_Sorter100|10414_ ;
  assign \new_Sorter100|10515_  = \new_Sorter100|10415_  & \new_Sorter100|10416_ ;
  assign \new_Sorter100|10516_  = \new_Sorter100|10415_  | \new_Sorter100|10416_ ;
  assign \new_Sorter100|10517_  = \new_Sorter100|10417_  & \new_Sorter100|10418_ ;
  assign \new_Sorter100|10518_  = \new_Sorter100|10417_  | \new_Sorter100|10418_ ;
  assign \new_Sorter100|10519_  = \new_Sorter100|10419_  & \new_Sorter100|10420_ ;
  assign \new_Sorter100|10520_  = \new_Sorter100|10419_  | \new_Sorter100|10420_ ;
  assign \new_Sorter100|10521_  = \new_Sorter100|10421_  & \new_Sorter100|10422_ ;
  assign \new_Sorter100|10522_  = \new_Sorter100|10421_  | \new_Sorter100|10422_ ;
  assign \new_Sorter100|10523_  = \new_Sorter100|10423_  & \new_Sorter100|10424_ ;
  assign \new_Sorter100|10524_  = \new_Sorter100|10423_  | \new_Sorter100|10424_ ;
  assign \new_Sorter100|10525_  = \new_Sorter100|10425_  & \new_Sorter100|10426_ ;
  assign \new_Sorter100|10526_  = \new_Sorter100|10425_  | \new_Sorter100|10426_ ;
  assign \new_Sorter100|10527_  = \new_Sorter100|10427_  & \new_Sorter100|10428_ ;
  assign \new_Sorter100|10528_  = \new_Sorter100|10427_  | \new_Sorter100|10428_ ;
  assign \new_Sorter100|10529_  = \new_Sorter100|10429_  & \new_Sorter100|10430_ ;
  assign \new_Sorter100|10530_  = \new_Sorter100|10429_  | \new_Sorter100|10430_ ;
  assign \new_Sorter100|10531_  = \new_Sorter100|10431_  & \new_Sorter100|10432_ ;
  assign \new_Sorter100|10532_  = \new_Sorter100|10431_  | \new_Sorter100|10432_ ;
  assign \new_Sorter100|10533_  = \new_Sorter100|10433_  & \new_Sorter100|10434_ ;
  assign \new_Sorter100|10534_  = \new_Sorter100|10433_  | \new_Sorter100|10434_ ;
  assign \new_Sorter100|10535_  = \new_Sorter100|10435_  & \new_Sorter100|10436_ ;
  assign \new_Sorter100|10536_  = \new_Sorter100|10435_  | \new_Sorter100|10436_ ;
  assign \new_Sorter100|10537_  = \new_Sorter100|10437_  & \new_Sorter100|10438_ ;
  assign \new_Sorter100|10538_  = \new_Sorter100|10437_  | \new_Sorter100|10438_ ;
  assign \new_Sorter100|10539_  = \new_Sorter100|10439_  & \new_Sorter100|10440_ ;
  assign \new_Sorter100|10540_  = \new_Sorter100|10439_  | \new_Sorter100|10440_ ;
  assign \new_Sorter100|10541_  = \new_Sorter100|10441_  & \new_Sorter100|10442_ ;
  assign \new_Sorter100|10542_  = \new_Sorter100|10441_  | \new_Sorter100|10442_ ;
  assign \new_Sorter100|10543_  = \new_Sorter100|10443_  & \new_Sorter100|10444_ ;
  assign \new_Sorter100|10544_  = \new_Sorter100|10443_  | \new_Sorter100|10444_ ;
  assign \new_Sorter100|10545_  = \new_Sorter100|10445_  & \new_Sorter100|10446_ ;
  assign \new_Sorter100|10546_  = \new_Sorter100|10445_  | \new_Sorter100|10446_ ;
  assign \new_Sorter100|10547_  = \new_Sorter100|10447_  & \new_Sorter100|10448_ ;
  assign \new_Sorter100|10548_  = \new_Sorter100|10447_  | \new_Sorter100|10448_ ;
  assign \new_Sorter100|10549_  = \new_Sorter100|10449_  & \new_Sorter100|10450_ ;
  assign \new_Sorter100|10550_  = \new_Sorter100|10449_  | \new_Sorter100|10450_ ;
  assign \new_Sorter100|10551_  = \new_Sorter100|10451_  & \new_Sorter100|10452_ ;
  assign \new_Sorter100|10552_  = \new_Sorter100|10451_  | \new_Sorter100|10452_ ;
  assign \new_Sorter100|10553_  = \new_Sorter100|10453_  & \new_Sorter100|10454_ ;
  assign \new_Sorter100|10554_  = \new_Sorter100|10453_  | \new_Sorter100|10454_ ;
  assign \new_Sorter100|10555_  = \new_Sorter100|10455_  & \new_Sorter100|10456_ ;
  assign \new_Sorter100|10556_  = \new_Sorter100|10455_  | \new_Sorter100|10456_ ;
  assign \new_Sorter100|10557_  = \new_Sorter100|10457_  & \new_Sorter100|10458_ ;
  assign \new_Sorter100|10558_  = \new_Sorter100|10457_  | \new_Sorter100|10458_ ;
  assign \new_Sorter100|10559_  = \new_Sorter100|10459_  & \new_Sorter100|10460_ ;
  assign \new_Sorter100|10560_  = \new_Sorter100|10459_  | \new_Sorter100|10460_ ;
  assign \new_Sorter100|10561_  = \new_Sorter100|10461_  & \new_Sorter100|10462_ ;
  assign \new_Sorter100|10562_  = \new_Sorter100|10461_  | \new_Sorter100|10462_ ;
  assign \new_Sorter100|10563_  = \new_Sorter100|10463_  & \new_Sorter100|10464_ ;
  assign \new_Sorter100|10564_  = \new_Sorter100|10463_  | \new_Sorter100|10464_ ;
  assign \new_Sorter100|10565_  = \new_Sorter100|10465_  & \new_Sorter100|10466_ ;
  assign \new_Sorter100|10566_  = \new_Sorter100|10465_  | \new_Sorter100|10466_ ;
  assign \new_Sorter100|10567_  = \new_Sorter100|10467_  & \new_Sorter100|10468_ ;
  assign \new_Sorter100|10568_  = \new_Sorter100|10467_  | \new_Sorter100|10468_ ;
  assign \new_Sorter100|10569_  = \new_Sorter100|10469_  & \new_Sorter100|10470_ ;
  assign \new_Sorter100|10570_  = \new_Sorter100|10469_  | \new_Sorter100|10470_ ;
  assign \new_Sorter100|10571_  = \new_Sorter100|10471_  & \new_Sorter100|10472_ ;
  assign \new_Sorter100|10572_  = \new_Sorter100|10471_  | \new_Sorter100|10472_ ;
  assign \new_Sorter100|10573_  = \new_Sorter100|10473_  & \new_Sorter100|10474_ ;
  assign \new_Sorter100|10574_  = \new_Sorter100|10473_  | \new_Sorter100|10474_ ;
  assign \new_Sorter100|10575_  = \new_Sorter100|10475_  & \new_Sorter100|10476_ ;
  assign \new_Sorter100|10576_  = \new_Sorter100|10475_  | \new_Sorter100|10476_ ;
  assign \new_Sorter100|10577_  = \new_Sorter100|10477_  & \new_Sorter100|10478_ ;
  assign \new_Sorter100|10578_  = \new_Sorter100|10477_  | \new_Sorter100|10478_ ;
  assign \new_Sorter100|10579_  = \new_Sorter100|10479_  & \new_Sorter100|10480_ ;
  assign \new_Sorter100|10580_  = \new_Sorter100|10479_  | \new_Sorter100|10480_ ;
  assign \new_Sorter100|10581_  = \new_Sorter100|10481_  & \new_Sorter100|10482_ ;
  assign \new_Sorter100|10582_  = \new_Sorter100|10481_  | \new_Sorter100|10482_ ;
  assign \new_Sorter100|10583_  = \new_Sorter100|10483_  & \new_Sorter100|10484_ ;
  assign \new_Sorter100|10584_  = \new_Sorter100|10483_  | \new_Sorter100|10484_ ;
  assign \new_Sorter100|10585_  = \new_Sorter100|10485_  & \new_Sorter100|10486_ ;
  assign \new_Sorter100|10586_  = \new_Sorter100|10485_  | \new_Sorter100|10486_ ;
  assign \new_Sorter100|10587_  = \new_Sorter100|10487_  & \new_Sorter100|10488_ ;
  assign \new_Sorter100|10588_  = \new_Sorter100|10487_  | \new_Sorter100|10488_ ;
  assign \new_Sorter100|10589_  = \new_Sorter100|10489_  & \new_Sorter100|10490_ ;
  assign \new_Sorter100|10590_  = \new_Sorter100|10489_  | \new_Sorter100|10490_ ;
  assign \new_Sorter100|10591_  = \new_Sorter100|10491_  & \new_Sorter100|10492_ ;
  assign \new_Sorter100|10592_  = \new_Sorter100|10491_  | \new_Sorter100|10492_ ;
  assign \new_Sorter100|10593_  = \new_Sorter100|10493_  & \new_Sorter100|10494_ ;
  assign \new_Sorter100|10594_  = \new_Sorter100|10493_  | \new_Sorter100|10494_ ;
  assign \new_Sorter100|10595_  = \new_Sorter100|10495_  & \new_Sorter100|10496_ ;
  assign \new_Sorter100|10596_  = \new_Sorter100|10495_  | \new_Sorter100|10496_ ;
  assign \new_Sorter100|10597_  = \new_Sorter100|10497_  & \new_Sorter100|10498_ ;
  assign \new_Sorter100|10598_  = \new_Sorter100|10497_  | \new_Sorter100|10498_ ;
  assign \new_Sorter100|10600_  = \new_Sorter100|10500_  & \new_Sorter100|10501_ ;
  assign \new_Sorter100|10601_  = \new_Sorter100|10500_  | \new_Sorter100|10501_ ;
  assign \new_Sorter100|10602_  = \new_Sorter100|10502_  & \new_Sorter100|10503_ ;
  assign \new_Sorter100|10603_  = \new_Sorter100|10502_  | \new_Sorter100|10503_ ;
  assign \new_Sorter100|10604_  = \new_Sorter100|10504_  & \new_Sorter100|10505_ ;
  assign \new_Sorter100|10605_  = \new_Sorter100|10504_  | \new_Sorter100|10505_ ;
  assign \new_Sorter100|10606_  = \new_Sorter100|10506_  & \new_Sorter100|10507_ ;
  assign \new_Sorter100|10607_  = \new_Sorter100|10506_  | \new_Sorter100|10507_ ;
  assign \new_Sorter100|10608_  = \new_Sorter100|10508_  & \new_Sorter100|10509_ ;
  assign \new_Sorter100|10609_  = \new_Sorter100|10508_  | \new_Sorter100|10509_ ;
  assign \new_Sorter100|10610_  = \new_Sorter100|10510_  & \new_Sorter100|10511_ ;
  assign \new_Sorter100|10611_  = \new_Sorter100|10510_  | \new_Sorter100|10511_ ;
  assign \new_Sorter100|10612_  = \new_Sorter100|10512_  & \new_Sorter100|10513_ ;
  assign \new_Sorter100|10613_  = \new_Sorter100|10512_  | \new_Sorter100|10513_ ;
  assign \new_Sorter100|10614_  = \new_Sorter100|10514_  & \new_Sorter100|10515_ ;
  assign \new_Sorter100|10615_  = \new_Sorter100|10514_  | \new_Sorter100|10515_ ;
  assign \new_Sorter100|10616_  = \new_Sorter100|10516_  & \new_Sorter100|10517_ ;
  assign \new_Sorter100|10617_  = \new_Sorter100|10516_  | \new_Sorter100|10517_ ;
  assign \new_Sorter100|10618_  = \new_Sorter100|10518_  & \new_Sorter100|10519_ ;
  assign \new_Sorter100|10619_  = \new_Sorter100|10518_  | \new_Sorter100|10519_ ;
  assign \new_Sorter100|10620_  = \new_Sorter100|10520_  & \new_Sorter100|10521_ ;
  assign \new_Sorter100|10621_  = \new_Sorter100|10520_  | \new_Sorter100|10521_ ;
  assign \new_Sorter100|10622_  = \new_Sorter100|10522_  & \new_Sorter100|10523_ ;
  assign \new_Sorter100|10623_  = \new_Sorter100|10522_  | \new_Sorter100|10523_ ;
  assign \new_Sorter100|10624_  = \new_Sorter100|10524_  & \new_Sorter100|10525_ ;
  assign \new_Sorter100|10625_  = \new_Sorter100|10524_  | \new_Sorter100|10525_ ;
  assign \new_Sorter100|10626_  = \new_Sorter100|10526_  & \new_Sorter100|10527_ ;
  assign \new_Sorter100|10627_  = \new_Sorter100|10526_  | \new_Sorter100|10527_ ;
  assign \new_Sorter100|10628_  = \new_Sorter100|10528_  & \new_Sorter100|10529_ ;
  assign \new_Sorter100|10629_  = \new_Sorter100|10528_  | \new_Sorter100|10529_ ;
  assign \new_Sorter100|10630_  = \new_Sorter100|10530_  & \new_Sorter100|10531_ ;
  assign \new_Sorter100|10631_  = \new_Sorter100|10530_  | \new_Sorter100|10531_ ;
  assign \new_Sorter100|10632_  = \new_Sorter100|10532_  & \new_Sorter100|10533_ ;
  assign \new_Sorter100|10633_  = \new_Sorter100|10532_  | \new_Sorter100|10533_ ;
  assign \new_Sorter100|10634_  = \new_Sorter100|10534_  & \new_Sorter100|10535_ ;
  assign \new_Sorter100|10635_  = \new_Sorter100|10534_  | \new_Sorter100|10535_ ;
  assign \new_Sorter100|10636_  = \new_Sorter100|10536_  & \new_Sorter100|10537_ ;
  assign \new_Sorter100|10637_  = \new_Sorter100|10536_  | \new_Sorter100|10537_ ;
  assign \new_Sorter100|10638_  = \new_Sorter100|10538_  & \new_Sorter100|10539_ ;
  assign \new_Sorter100|10639_  = \new_Sorter100|10538_  | \new_Sorter100|10539_ ;
  assign \new_Sorter100|10640_  = \new_Sorter100|10540_  & \new_Sorter100|10541_ ;
  assign \new_Sorter100|10641_  = \new_Sorter100|10540_  | \new_Sorter100|10541_ ;
  assign \new_Sorter100|10642_  = \new_Sorter100|10542_  & \new_Sorter100|10543_ ;
  assign \new_Sorter100|10643_  = \new_Sorter100|10542_  | \new_Sorter100|10543_ ;
  assign \new_Sorter100|10644_  = \new_Sorter100|10544_  & \new_Sorter100|10545_ ;
  assign \new_Sorter100|10645_  = \new_Sorter100|10544_  | \new_Sorter100|10545_ ;
  assign \new_Sorter100|10646_  = \new_Sorter100|10546_  & \new_Sorter100|10547_ ;
  assign \new_Sorter100|10647_  = \new_Sorter100|10546_  | \new_Sorter100|10547_ ;
  assign \new_Sorter100|10648_  = \new_Sorter100|10548_  & \new_Sorter100|10549_ ;
  assign \new_Sorter100|10649_  = \new_Sorter100|10548_  | \new_Sorter100|10549_ ;
  assign \new_Sorter100|10650_  = \new_Sorter100|10550_  & \new_Sorter100|10551_ ;
  assign \new_Sorter100|10651_  = \new_Sorter100|10550_  | \new_Sorter100|10551_ ;
  assign \new_Sorter100|10652_  = \new_Sorter100|10552_  & \new_Sorter100|10553_ ;
  assign \new_Sorter100|10653_  = \new_Sorter100|10552_  | \new_Sorter100|10553_ ;
  assign \new_Sorter100|10654_  = \new_Sorter100|10554_  & \new_Sorter100|10555_ ;
  assign \new_Sorter100|10655_  = \new_Sorter100|10554_  | \new_Sorter100|10555_ ;
  assign \new_Sorter100|10656_  = \new_Sorter100|10556_  & \new_Sorter100|10557_ ;
  assign \new_Sorter100|10657_  = \new_Sorter100|10556_  | \new_Sorter100|10557_ ;
  assign \new_Sorter100|10658_  = \new_Sorter100|10558_  & \new_Sorter100|10559_ ;
  assign \new_Sorter100|10659_  = \new_Sorter100|10558_  | \new_Sorter100|10559_ ;
  assign \new_Sorter100|10660_  = \new_Sorter100|10560_  & \new_Sorter100|10561_ ;
  assign \new_Sorter100|10661_  = \new_Sorter100|10560_  | \new_Sorter100|10561_ ;
  assign \new_Sorter100|10662_  = \new_Sorter100|10562_  & \new_Sorter100|10563_ ;
  assign \new_Sorter100|10663_  = \new_Sorter100|10562_  | \new_Sorter100|10563_ ;
  assign \new_Sorter100|10664_  = \new_Sorter100|10564_  & \new_Sorter100|10565_ ;
  assign \new_Sorter100|10665_  = \new_Sorter100|10564_  | \new_Sorter100|10565_ ;
  assign \new_Sorter100|10666_  = \new_Sorter100|10566_  & \new_Sorter100|10567_ ;
  assign \new_Sorter100|10667_  = \new_Sorter100|10566_  | \new_Sorter100|10567_ ;
  assign \new_Sorter100|10668_  = \new_Sorter100|10568_  & \new_Sorter100|10569_ ;
  assign \new_Sorter100|10669_  = \new_Sorter100|10568_  | \new_Sorter100|10569_ ;
  assign \new_Sorter100|10670_  = \new_Sorter100|10570_  & \new_Sorter100|10571_ ;
  assign \new_Sorter100|10671_  = \new_Sorter100|10570_  | \new_Sorter100|10571_ ;
  assign \new_Sorter100|10672_  = \new_Sorter100|10572_  & \new_Sorter100|10573_ ;
  assign \new_Sorter100|10673_  = \new_Sorter100|10572_  | \new_Sorter100|10573_ ;
  assign \new_Sorter100|10674_  = \new_Sorter100|10574_  & \new_Sorter100|10575_ ;
  assign \new_Sorter100|10675_  = \new_Sorter100|10574_  | \new_Sorter100|10575_ ;
  assign \new_Sorter100|10676_  = \new_Sorter100|10576_  & \new_Sorter100|10577_ ;
  assign \new_Sorter100|10677_  = \new_Sorter100|10576_  | \new_Sorter100|10577_ ;
  assign \new_Sorter100|10678_  = \new_Sorter100|10578_  & \new_Sorter100|10579_ ;
  assign \new_Sorter100|10679_  = \new_Sorter100|10578_  | \new_Sorter100|10579_ ;
  assign \new_Sorter100|10680_  = \new_Sorter100|10580_  & \new_Sorter100|10581_ ;
  assign \new_Sorter100|10681_  = \new_Sorter100|10580_  | \new_Sorter100|10581_ ;
  assign \new_Sorter100|10682_  = \new_Sorter100|10582_  & \new_Sorter100|10583_ ;
  assign \new_Sorter100|10683_  = \new_Sorter100|10582_  | \new_Sorter100|10583_ ;
  assign \new_Sorter100|10684_  = \new_Sorter100|10584_  & \new_Sorter100|10585_ ;
  assign \new_Sorter100|10685_  = \new_Sorter100|10584_  | \new_Sorter100|10585_ ;
  assign \new_Sorter100|10686_  = \new_Sorter100|10586_  & \new_Sorter100|10587_ ;
  assign \new_Sorter100|10687_  = \new_Sorter100|10586_  | \new_Sorter100|10587_ ;
  assign \new_Sorter100|10688_  = \new_Sorter100|10588_  & \new_Sorter100|10589_ ;
  assign \new_Sorter100|10689_  = \new_Sorter100|10588_  | \new_Sorter100|10589_ ;
  assign \new_Sorter100|10690_  = \new_Sorter100|10590_  & \new_Sorter100|10591_ ;
  assign \new_Sorter100|10691_  = \new_Sorter100|10590_  | \new_Sorter100|10591_ ;
  assign \new_Sorter100|10692_  = \new_Sorter100|10592_  & \new_Sorter100|10593_ ;
  assign \new_Sorter100|10693_  = \new_Sorter100|10592_  | \new_Sorter100|10593_ ;
  assign \new_Sorter100|10694_  = \new_Sorter100|10594_  & \new_Sorter100|10595_ ;
  assign \new_Sorter100|10695_  = \new_Sorter100|10594_  | \new_Sorter100|10595_ ;
  assign \new_Sorter100|10696_  = \new_Sorter100|10596_  & \new_Sorter100|10597_ ;
  assign \new_Sorter100|10697_  = \new_Sorter100|10596_  | \new_Sorter100|10597_ ;
  assign \new_Sorter100|10698_  = \new_Sorter100|10598_  & \new_Sorter100|10599_ ;
  assign \new_Sorter100|10699_  = \new_Sorter100|10598_  | \new_Sorter100|10599_ ;
  assign \new_Sorter100|10700_  = \new_Sorter100|10600_ ;
  assign \new_Sorter100|10799_  = \new_Sorter100|10699_ ;
  assign \new_Sorter100|10701_  = \new_Sorter100|10601_  & \new_Sorter100|10602_ ;
  assign \new_Sorter100|10702_  = \new_Sorter100|10601_  | \new_Sorter100|10602_ ;
  assign \new_Sorter100|10703_  = \new_Sorter100|10603_  & \new_Sorter100|10604_ ;
  assign \new_Sorter100|10704_  = \new_Sorter100|10603_  | \new_Sorter100|10604_ ;
  assign \new_Sorter100|10705_  = \new_Sorter100|10605_  & \new_Sorter100|10606_ ;
  assign \new_Sorter100|10706_  = \new_Sorter100|10605_  | \new_Sorter100|10606_ ;
  assign \new_Sorter100|10707_  = \new_Sorter100|10607_  & \new_Sorter100|10608_ ;
  assign \new_Sorter100|10708_  = \new_Sorter100|10607_  | \new_Sorter100|10608_ ;
  assign \new_Sorter100|10709_  = \new_Sorter100|10609_  & \new_Sorter100|10610_ ;
  assign \new_Sorter100|10710_  = \new_Sorter100|10609_  | \new_Sorter100|10610_ ;
  assign \new_Sorter100|10711_  = \new_Sorter100|10611_  & \new_Sorter100|10612_ ;
  assign \new_Sorter100|10712_  = \new_Sorter100|10611_  | \new_Sorter100|10612_ ;
  assign \new_Sorter100|10713_  = \new_Sorter100|10613_  & \new_Sorter100|10614_ ;
  assign \new_Sorter100|10714_  = \new_Sorter100|10613_  | \new_Sorter100|10614_ ;
  assign \new_Sorter100|10715_  = \new_Sorter100|10615_  & \new_Sorter100|10616_ ;
  assign \new_Sorter100|10716_  = \new_Sorter100|10615_  | \new_Sorter100|10616_ ;
  assign \new_Sorter100|10717_  = \new_Sorter100|10617_  & \new_Sorter100|10618_ ;
  assign \new_Sorter100|10718_  = \new_Sorter100|10617_  | \new_Sorter100|10618_ ;
  assign \new_Sorter100|10719_  = \new_Sorter100|10619_  & \new_Sorter100|10620_ ;
  assign \new_Sorter100|10720_  = \new_Sorter100|10619_  | \new_Sorter100|10620_ ;
  assign \new_Sorter100|10721_  = \new_Sorter100|10621_  & \new_Sorter100|10622_ ;
  assign \new_Sorter100|10722_  = \new_Sorter100|10621_  | \new_Sorter100|10622_ ;
  assign \new_Sorter100|10723_  = \new_Sorter100|10623_  & \new_Sorter100|10624_ ;
  assign \new_Sorter100|10724_  = \new_Sorter100|10623_  | \new_Sorter100|10624_ ;
  assign \new_Sorter100|10725_  = \new_Sorter100|10625_  & \new_Sorter100|10626_ ;
  assign \new_Sorter100|10726_  = \new_Sorter100|10625_  | \new_Sorter100|10626_ ;
  assign \new_Sorter100|10727_  = \new_Sorter100|10627_  & \new_Sorter100|10628_ ;
  assign \new_Sorter100|10728_  = \new_Sorter100|10627_  | \new_Sorter100|10628_ ;
  assign \new_Sorter100|10729_  = \new_Sorter100|10629_  & \new_Sorter100|10630_ ;
  assign \new_Sorter100|10730_  = \new_Sorter100|10629_  | \new_Sorter100|10630_ ;
  assign \new_Sorter100|10731_  = \new_Sorter100|10631_  & \new_Sorter100|10632_ ;
  assign \new_Sorter100|10732_  = \new_Sorter100|10631_  | \new_Sorter100|10632_ ;
  assign \new_Sorter100|10733_  = \new_Sorter100|10633_  & \new_Sorter100|10634_ ;
  assign \new_Sorter100|10734_  = \new_Sorter100|10633_  | \new_Sorter100|10634_ ;
  assign \new_Sorter100|10735_  = \new_Sorter100|10635_  & \new_Sorter100|10636_ ;
  assign \new_Sorter100|10736_  = \new_Sorter100|10635_  | \new_Sorter100|10636_ ;
  assign \new_Sorter100|10737_  = \new_Sorter100|10637_  & \new_Sorter100|10638_ ;
  assign \new_Sorter100|10738_  = \new_Sorter100|10637_  | \new_Sorter100|10638_ ;
  assign \new_Sorter100|10739_  = \new_Sorter100|10639_  & \new_Sorter100|10640_ ;
  assign \new_Sorter100|10740_  = \new_Sorter100|10639_  | \new_Sorter100|10640_ ;
  assign \new_Sorter100|10741_  = \new_Sorter100|10641_  & \new_Sorter100|10642_ ;
  assign \new_Sorter100|10742_  = \new_Sorter100|10641_  | \new_Sorter100|10642_ ;
  assign \new_Sorter100|10743_  = \new_Sorter100|10643_  & \new_Sorter100|10644_ ;
  assign \new_Sorter100|10744_  = \new_Sorter100|10643_  | \new_Sorter100|10644_ ;
  assign \new_Sorter100|10745_  = \new_Sorter100|10645_  & \new_Sorter100|10646_ ;
  assign \new_Sorter100|10746_  = \new_Sorter100|10645_  | \new_Sorter100|10646_ ;
  assign \new_Sorter100|10747_  = \new_Sorter100|10647_  & \new_Sorter100|10648_ ;
  assign \new_Sorter100|10748_  = \new_Sorter100|10647_  | \new_Sorter100|10648_ ;
  assign \new_Sorter100|10749_  = \new_Sorter100|10649_  & \new_Sorter100|10650_ ;
  assign \new_Sorter100|10750_  = \new_Sorter100|10649_  | \new_Sorter100|10650_ ;
  assign \new_Sorter100|10751_  = \new_Sorter100|10651_  & \new_Sorter100|10652_ ;
  assign \new_Sorter100|10752_  = \new_Sorter100|10651_  | \new_Sorter100|10652_ ;
  assign \new_Sorter100|10753_  = \new_Sorter100|10653_  & \new_Sorter100|10654_ ;
  assign \new_Sorter100|10754_  = \new_Sorter100|10653_  | \new_Sorter100|10654_ ;
  assign \new_Sorter100|10755_  = \new_Sorter100|10655_  & \new_Sorter100|10656_ ;
  assign \new_Sorter100|10756_  = \new_Sorter100|10655_  | \new_Sorter100|10656_ ;
  assign \new_Sorter100|10757_  = \new_Sorter100|10657_  & \new_Sorter100|10658_ ;
  assign \new_Sorter100|10758_  = \new_Sorter100|10657_  | \new_Sorter100|10658_ ;
  assign \new_Sorter100|10759_  = \new_Sorter100|10659_  & \new_Sorter100|10660_ ;
  assign \new_Sorter100|10760_  = \new_Sorter100|10659_  | \new_Sorter100|10660_ ;
  assign \new_Sorter100|10761_  = \new_Sorter100|10661_  & \new_Sorter100|10662_ ;
  assign \new_Sorter100|10762_  = \new_Sorter100|10661_  | \new_Sorter100|10662_ ;
  assign \new_Sorter100|10763_  = \new_Sorter100|10663_  & \new_Sorter100|10664_ ;
  assign \new_Sorter100|10764_  = \new_Sorter100|10663_  | \new_Sorter100|10664_ ;
  assign \new_Sorter100|10765_  = \new_Sorter100|10665_  & \new_Sorter100|10666_ ;
  assign \new_Sorter100|10766_  = \new_Sorter100|10665_  | \new_Sorter100|10666_ ;
  assign \new_Sorter100|10767_  = \new_Sorter100|10667_  & \new_Sorter100|10668_ ;
  assign \new_Sorter100|10768_  = \new_Sorter100|10667_  | \new_Sorter100|10668_ ;
  assign \new_Sorter100|10769_  = \new_Sorter100|10669_  & \new_Sorter100|10670_ ;
  assign \new_Sorter100|10770_  = \new_Sorter100|10669_  | \new_Sorter100|10670_ ;
  assign \new_Sorter100|10771_  = \new_Sorter100|10671_  & \new_Sorter100|10672_ ;
  assign \new_Sorter100|10772_  = \new_Sorter100|10671_  | \new_Sorter100|10672_ ;
  assign \new_Sorter100|10773_  = \new_Sorter100|10673_  & \new_Sorter100|10674_ ;
  assign \new_Sorter100|10774_  = \new_Sorter100|10673_  | \new_Sorter100|10674_ ;
  assign \new_Sorter100|10775_  = \new_Sorter100|10675_  & \new_Sorter100|10676_ ;
  assign \new_Sorter100|10776_  = \new_Sorter100|10675_  | \new_Sorter100|10676_ ;
  assign \new_Sorter100|10777_  = \new_Sorter100|10677_  & \new_Sorter100|10678_ ;
  assign \new_Sorter100|10778_  = \new_Sorter100|10677_  | \new_Sorter100|10678_ ;
  assign \new_Sorter100|10779_  = \new_Sorter100|10679_  & \new_Sorter100|10680_ ;
  assign \new_Sorter100|10780_  = \new_Sorter100|10679_  | \new_Sorter100|10680_ ;
  assign \new_Sorter100|10781_  = \new_Sorter100|10681_  & \new_Sorter100|10682_ ;
  assign \new_Sorter100|10782_  = \new_Sorter100|10681_  | \new_Sorter100|10682_ ;
  assign \new_Sorter100|10783_  = \new_Sorter100|10683_  & \new_Sorter100|10684_ ;
  assign \new_Sorter100|10784_  = \new_Sorter100|10683_  | \new_Sorter100|10684_ ;
  assign \new_Sorter100|10785_  = \new_Sorter100|10685_  & \new_Sorter100|10686_ ;
  assign \new_Sorter100|10786_  = \new_Sorter100|10685_  | \new_Sorter100|10686_ ;
  assign \new_Sorter100|10787_  = \new_Sorter100|10687_  & \new_Sorter100|10688_ ;
  assign \new_Sorter100|10788_  = \new_Sorter100|10687_  | \new_Sorter100|10688_ ;
  assign \new_Sorter100|10789_  = \new_Sorter100|10689_  & \new_Sorter100|10690_ ;
  assign \new_Sorter100|10790_  = \new_Sorter100|10689_  | \new_Sorter100|10690_ ;
  assign \new_Sorter100|10791_  = \new_Sorter100|10691_  & \new_Sorter100|10692_ ;
  assign \new_Sorter100|10792_  = \new_Sorter100|10691_  | \new_Sorter100|10692_ ;
  assign \new_Sorter100|10793_  = \new_Sorter100|10693_  & \new_Sorter100|10694_ ;
  assign \new_Sorter100|10794_  = \new_Sorter100|10693_  | \new_Sorter100|10694_ ;
  assign \new_Sorter100|10795_  = \new_Sorter100|10695_  & \new_Sorter100|10696_ ;
  assign \new_Sorter100|10796_  = \new_Sorter100|10695_  | \new_Sorter100|10696_ ;
  assign \new_Sorter100|10797_  = \new_Sorter100|10697_  & \new_Sorter100|10698_ ;
  assign \new_Sorter100|10798_  = \new_Sorter100|10697_  | \new_Sorter100|10698_ ;
  assign \new_Sorter100|10800_  = \new_Sorter100|10700_  & \new_Sorter100|10701_ ;
  assign \new_Sorter100|10801_  = \new_Sorter100|10700_  | \new_Sorter100|10701_ ;
  assign \new_Sorter100|10802_  = \new_Sorter100|10702_  & \new_Sorter100|10703_ ;
  assign \new_Sorter100|10803_  = \new_Sorter100|10702_  | \new_Sorter100|10703_ ;
  assign \new_Sorter100|10804_  = \new_Sorter100|10704_  & \new_Sorter100|10705_ ;
  assign \new_Sorter100|10805_  = \new_Sorter100|10704_  | \new_Sorter100|10705_ ;
  assign \new_Sorter100|10806_  = \new_Sorter100|10706_  & \new_Sorter100|10707_ ;
  assign \new_Sorter100|10807_  = \new_Sorter100|10706_  | \new_Sorter100|10707_ ;
  assign \new_Sorter100|10808_  = \new_Sorter100|10708_  & \new_Sorter100|10709_ ;
  assign \new_Sorter100|10809_  = \new_Sorter100|10708_  | \new_Sorter100|10709_ ;
  assign \new_Sorter100|10810_  = \new_Sorter100|10710_  & \new_Sorter100|10711_ ;
  assign \new_Sorter100|10811_  = \new_Sorter100|10710_  | \new_Sorter100|10711_ ;
  assign \new_Sorter100|10812_  = \new_Sorter100|10712_  & \new_Sorter100|10713_ ;
  assign \new_Sorter100|10813_  = \new_Sorter100|10712_  | \new_Sorter100|10713_ ;
  assign \new_Sorter100|10814_  = \new_Sorter100|10714_  & \new_Sorter100|10715_ ;
  assign \new_Sorter100|10815_  = \new_Sorter100|10714_  | \new_Sorter100|10715_ ;
  assign \new_Sorter100|10816_  = \new_Sorter100|10716_  & \new_Sorter100|10717_ ;
  assign \new_Sorter100|10817_  = \new_Sorter100|10716_  | \new_Sorter100|10717_ ;
  assign \new_Sorter100|10818_  = \new_Sorter100|10718_  & \new_Sorter100|10719_ ;
  assign \new_Sorter100|10819_  = \new_Sorter100|10718_  | \new_Sorter100|10719_ ;
  assign \new_Sorter100|10820_  = \new_Sorter100|10720_  & \new_Sorter100|10721_ ;
  assign \new_Sorter100|10821_  = \new_Sorter100|10720_  | \new_Sorter100|10721_ ;
  assign \new_Sorter100|10822_  = \new_Sorter100|10722_  & \new_Sorter100|10723_ ;
  assign \new_Sorter100|10823_  = \new_Sorter100|10722_  | \new_Sorter100|10723_ ;
  assign \new_Sorter100|10824_  = \new_Sorter100|10724_  & \new_Sorter100|10725_ ;
  assign \new_Sorter100|10825_  = \new_Sorter100|10724_  | \new_Sorter100|10725_ ;
  assign \new_Sorter100|10826_  = \new_Sorter100|10726_  & \new_Sorter100|10727_ ;
  assign \new_Sorter100|10827_  = \new_Sorter100|10726_  | \new_Sorter100|10727_ ;
  assign \new_Sorter100|10828_  = \new_Sorter100|10728_  & \new_Sorter100|10729_ ;
  assign \new_Sorter100|10829_  = \new_Sorter100|10728_  | \new_Sorter100|10729_ ;
  assign \new_Sorter100|10830_  = \new_Sorter100|10730_  & \new_Sorter100|10731_ ;
  assign \new_Sorter100|10831_  = \new_Sorter100|10730_  | \new_Sorter100|10731_ ;
  assign \new_Sorter100|10832_  = \new_Sorter100|10732_  & \new_Sorter100|10733_ ;
  assign \new_Sorter100|10833_  = \new_Sorter100|10732_  | \new_Sorter100|10733_ ;
  assign \new_Sorter100|10834_  = \new_Sorter100|10734_  & \new_Sorter100|10735_ ;
  assign \new_Sorter100|10835_  = \new_Sorter100|10734_  | \new_Sorter100|10735_ ;
  assign \new_Sorter100|10836_  = \new_Sorter100|10736_  & \new_Sorter100|10737_ ;
  assign \new_Sorter100|10837_  = \new_Sorter100|10736_  | \new_Sorter100|10737_ ;
  assign \new_Sorter100|10838_  = \new_Sorter100|10738_  & \new_Sorter100|10739_ ;
  assign \new_Sorter100|10839_  = \new_Sorter100|10738_  | \new_Sorter100|10739_ ;
  assign \new_Sorter100|10840_  = \new_Sorter100|10740_  & \new_Sorter100|10741_ ;
  assign \new_Sorter100|10841_  = \new_Sorter100|10740_  | \new_Sorter100|10741_ ;
  assign \new_Sorter100|10842_  = \new_Sorter100|10742_  & \new_Sorter100|10743_ ;
  assign \new_Sorter100|10843_  = \new_Sorter100|10742_  | \new_Sorter100|10743_ ;
  assign \new_Sorter100|10844_  = \new_Sorter100|10744_  & \new_Sorter100|10745_ ;
  assign \new_Sorter100|10845_  = \new_Sorter100|10744_  | \new_Sorter100|10745_ ;
  assign \new_Sorter100|10846_  = \new_Sorter100|10746_  & \new_Sorter100|10747_ ;
  assign \new_Sorter100|10847_  = \new_Sorter100|10746_  | \new_Sorter100|10747_ ;
  assign \new_Sorter100|10848_  = \new_Sorter100|10748_  & \new_Sorter100|10749_ ;
  assign \new_Sorter100|10849_  = \new_Sorter100|10748_  | \new_Sorter100|10749_ ;
  assign \new_Sorter100|10850_  = \new_Sorter100|10750_  & \new_Sorter100|10751_ ;
  assign \new_Sorter100|10851_  = \new_Sorter100|10750_  | \new_Sorter100|10751_ ;
  assign \new_Sorter100|10852_  = \new_Sorter100|10752_  & \new_Sorter100|10753_ ;
  assign \new_Sorter100|10853_  = \new_Sorter100|10752_  | \new_Sorter100|10753_ ;
  assign \new_Sorter100|10854_  = \new_Sorter100|10754_  & \new_Sorter100|10755_ ;
  assign \new_Sorter100|10855_  = \new_Sorter100|10754_  | \new_Sorter100|10755_ ;
  assign \new_Sorter100|10856_  = \new_Sorter100|10756_  & \new_Sorter100|10757_ ;
  assign \new_Sorter100|10857_  = \new_Sorter100|10756_  | \new_Sorter100|10757_ ;
  assign \new_Sorter100|10858_  = \new_Sorter100|10758_  & \new_Sorter100|10759_ ;
  assign \new_Sorter100|10859_  = \new_Sorter100|10758_  | \new_Sorter100|10759_ ;
  assign \new_Sorter100|10860_  = \new_Sorter100|10760_  & \new_Sorter100|10761_ ;
  assign \new_Sorter100|10861_  = \new_Sorter100|10760_  | \new_Sorter100|10761_ ;
  assign \new_Sorter100|10862_  = \new_Sorter100|10762_  & \new_Sorter100|10763_ ;
  assign \new_Sorter100|10863_  = \new_Sorter100|10762_  | \new_Sorter100|10763_ ;
  assign \new_Sorter100|10864_  = \new_Sorter100|10764_  & \new_Sorter100|10765_ ;
  assign \new_Sorter100|10865_  = \new_Sorter100|10764_  | \new_Sorter100|10765_ ;
  assign \new_Sorter100|10866_  = \new_Sorter100|10766_  & \new_Sorter100|10767_ ;
  assign \new_Sorter100|10867_  = \new_Sorter100|10766_  | \new_Sorter100|10767_ ;
  assign \new_Sorter100|10868_  = \new_Sorter100|10768_  & \new_Sorter100|10769_ ;
  assign \new_Sorter100|10869_  = \new_Sorter100|10768_  | \new_Sorter100|10769_ ;
  assign \new_Sorter100|10870_  = \new_Sorter100|10770_  & \new_Sorter100|10771_ ;
  assign \new_Sorter100|10871_  = \new_Sorter100|10770_  | \new_Sorter100|10771_ ;
  assign \new_Sorter100|10872_  = \new_Sorter100|10772_  & \new_Sorter100|10773_ ;
  assign \new_Sorter100|10873_  = \new_Sorter100|10772_  | \new_Sorter100|10773_ ;
  assign \new_Sorter100|10874_  = \new_Sorter100|10774_  & \new_Sorter100|10775_ ;
  assign \new_Sorter100|10875_  = \new_Sorter100|10774_  | \new_Sorter100|10775_ ;
  assign \new_Sorter100|10876_  = \new_Sorter100|10776_  & \new_Sorter100|10777_ ;
  assign \new_Sorter100|10877_  = \new_Sorter100|10776_  | \new_Sorter100|10777_ ;
  assign \new_Sorter100|10878_  = \new_Sorter100|10778_  & \new_Sorter100|10779_ ;
  assign \new_Sorter100|10879_  = \new_Sorter100|10778_  | \new_Sorter100|10779_ ;
  assign \new_Sorter100|10880_  = \new_Sorter100|10780_  & \new_Sorter100|10781_ ;
  assign \new_Sorter100|10881_  = \new_Sorter100|10780_  | \new_Sorter100|10781_ ;
  assign \new_Sorter100|10882_  = \new_Sorter100|10782_  & \new_Sorter100|10783_ ;
  assign \new_Sorter100|10883_  = \new_Sorter100|10782_  | \new_Sorter100|10783_ ;
  assign \new_Sorter100|10884_  = \new_Sorter100|10784_  & \new_Sorter100|10785_ ;
  assign \new_Sorter100|10885_  = \new_Sorter100|10784_  | \new_Sorter100|10785_ ;
  assign \new_Sorter100|10886_  = \new_Sorter100|10786_  & \new_Sorter100|10787_ ;
  assign \new_Sorter100|10887_  = \new_Sorter100|10786_  | \new_Sorter100|10787_ ;
  assign \new_Sorter100|10888_  = \new_Sorter100|10788_  & \new_Sorter100|10789_ ;
  assign \new_Sorter100|10889_  = \new_Sorter100|10788_  | \new_Sorter100|10789_ ;
  assign \new_Sorter100|10890_  = \new_Sorter100|10790_  & \new_Sorter100|10791_ ;
  assign \new_Sorter100|10891_  = \new_Sorter100|10790_  | \new_Sorter100|10791_ ;
  assign \new_Sorter100|10892_  = \new_Sorter100|10792_  & \new_Sorter100|10793_ ;
  assign \new_Sorter100|10893_  = \new_Sorter100|10792_  | \new_Sorter100|10793_ ;
  assign \new_Sorter100|10894_  = \new_Sorter100|10794_  & \new_Sorter100|10795_ ;
  assign \new_Sorter100|10895_  = \new_Sorter100|10794_  | \new_Sorter100|10795_ ;
  assign \new_Sorter100|10896_  = \new_Sorter100|10796_  & \new_Sorter100|10797_ ;
  assign \new_Sorter100|10897_  = \new_Sorter100|10796_  | \new_Sorter100|10797_ ;
  assign \new_Sorter100|10898_  = \new_Sorter100|10798_  & \new_Sorter100|10799_ ;
  assign \new_Sorter100|10899_  = \new_Sorter100|10798_  | \new_Sorter100|10799_ ;
  assign \new_Sorter100|10900_  = \new_Sorter100|10800_ ;
  assign \new_Sorter100|10999_  = \new_Sorter100|10899_ ;
  assign \new_Sorter100|10901_  = \new_Sorter100|10801_  & \new_Sorter100|10802_ ;
  assign \new_Sorter100|10902_  = \new_Sorter100|10801_  | \new_Sorter100|10802_ ;
  assign \new_Sorter100|10903_  = \new_Sorter100|10803_  & \new_Sorter100|10804_ ;
  assign \new_Sorter100|10904_  = \new_Sorter100|10803_  | \new_Sorter100|10804_ ;
  assign \new_Sorter100|10905_  = \new_Sorter100|10805_  & \new_Sorter100|10806_ ;
  assign \new_Sorter100|10906_  = \new_Sorter100|10805_  | \new_Sorter100|10806_ ;
  assign \new_Sorter100|10907_  = \new_Sorter100|10807_  & \new_Sorter100|10808_ ;
  assign \new_Sorter100|10908_  = \new_Sorter100|10807_  | \new_Sorter100|10808_ ;
  assign \new_Sorter100|10909_  = \new_Sorter100|10809_  & \new_Sorter100|10810_ ;
  assign \new_Sorter100|10910_  = \new_Sorter100|10809_  | \new_Sorter100|10810_ ;
  assign \new_Sorter100|10911_  = \new_Sorter100|10811_  & \new_Sorter100|10812_ ;
  assign \new_Sorter100|10912_  = \new_Sorter100|10811_  | \new_Sorter100|10812_ ;
  assign \new_Sorter100|10913_  = \new_Sorter100|10813_  & \new_Sorter100|10814_ ;
  assign \new_Sorter100|10914_  = \new_Sorter100|10813_  | \new_Sorter100|10814_ ;
  assign \new_Sorter100|10915_  = \new_Sorter100|10815_  & \new_Sorter100|10816_ ;
  assign \new_Sorter100|10916_  = \new_Sorter100|10815_  | \new_Sorter100|10816_ ;
  assign \new_Sorter100|10917_  = \new_Sorter100|10817_  & \new_Sorter100|10818_ ;
  assign \new_Sorter100|10918_  = \new_Sorter100|10817_  | \new_Sorter100|10818_ ;
  assign \new_Sorter100|10919_  = \new_Sorter100|10819_  & \new_Sorter100|10820_ ;
  assign \new_Sorter100|10920_  = \new_Sorter100|10819_  | \new_Sorter100|10820_ ;
  assign \new_Sorter100|10921_  = \new_Sorter100|10821_  & \new_Sorter100|10822_ ;
  assign \new_Sorter100|10922_  = \new_Sorter100|10821_  | \new_Sorter100|10822_ ;
  assign \new_Sorter100|10923_  = \new_Sorter100|10823_  & \new_Sorter100|10824_ ;
  assign \new_Sorter100|10924_  = \new_Sorter100|10823_  | \new_Sorter100|10824_ ;
  assign \new_Sorter100|10925_  = \new_Sorter100|10825_  & \new_Sorter100|10826_ ;
  assign \new_Sorter100|10926_  = \new_Sorter100|10825_  | \new_Sorter100|10826_ ;
  assign \new_Sorter100|10927_  = \new_Sorter100|10827_  & \new_Sorter100|10828_ ;
  assign \new_Sorter100|10928_  = \new_Sorter100|10827_  | \new_Sorter100|10828_ ;
  assign \new_Sorter100|10929_  = \new_Sorter100|10829_  & \new_Sorter100|10830_ ;
  assign \new_Sorter100|10930_  = \new_Sorter100|10829_  | \new_Sorter100|10830_ ;
  assign \new_Sorter100|10931_  = \new_Sorter100|10831_  & \new_Sorter100|10832_ ;
  assign \new_Sorter100|10932_  = \new_Sorter100|10831_  | \new_Sorter100|10832_ ;
  assign \new_Sorter100|10933_  = \new_Sorter100|10833_  & \new_Sorter100|10834_ ;
  assign \new_Sorter100|10934_  = \new_Sorter100|10833_  | \new_Sorter100|10834_ ;
  assign \new_Sorter100|10935_  = \new_Sorter100|10835_  & \new_Sorter100|10836_ ;
  assign \new_Sorter100|10936_  = \new_Sorter100|10835_  | \new_Sorter100|10836_ ;
  assign \new_Sorter100|10937_  = \new_Sorter100|10837_  & \new_Sorter100|10838_ ;
  assign \new_Sorter100|10938_  = \new_Sorter100|10837_  | \new_Sorter100|10838_ ;
  assign \new_Sorter100|10939_  = \new_Sorter100|10839_  & \new_Sorter100|10840_ ;
  assign \new_Sorter100|10940_  = \new_Sorter100|10839_  | \new_Sorter100|10840_ ;
  assign \new_Sorter100|10941_  = \new_Sorter100|10841_  & \new_Sorter100|10842_ ;
  assign \new_Sorter100|10942_  = \new_Sorter100|10841_  | \new_Sorter100|10842_ ;
  assign \new_Sorter100|10943_  = \new_Sorter100|10843_  & \new_Sorter100|10844_ ;
  assign \new_Sorter100|10944_  = \new_Sorter100|10843_  | \new_Sorter100|10844_ ;
  assign \new_Sorter100|10945_  = \new_Sorter100|10845_  & \new_Sorter100|10846_ ;
  assign \new_Sorter100|10946_  = \new_Sorter100|10845_  | \new_Sorter100|10846_ ;
  assign \new_Sorter100|10947_  = \new_Sorter100|10847_  & \new_Sorter100|10848_ ;
  assign \new_Sorter100|10948_  = \new_Sorter100|10847_  | \new_Sorter100|10848_ ;
  assign \new_Sorter100|10949_  = \new_Sorter100|10849_  & \new_Sorter100|10850_ ;
  assign \new_Sorter100|10950_  = \new_Sorter100|10849_  | \new_Sorter100|10850_ ;
  assign \new_Sorter100|10951_  = \new_Sorter100|10851_  & \new_Sorter100|10852_ ;
  assign \new_Sorter100|10952_  = \new_Sorter100|10851_  | \new_Sorter100|10852_ ;
  assign \new_Sorter100|10953_  = \new_Sorter100|10853_  & \new_Sorter100|10854_ ;
  assign \new_Sorter100|10954_  = \new_Sorter100|10853_  | \new_Sorter100|10854_ ;
  assign \new_Sorter100|10955_  = \new_Sorter100|10855_  & \new_Sorter100|10856_ ;
  assign \new_Sorter100|10956_  = \new_Sorter100|10855_  | \new_Sorter100|10856_ ;
  assign \new_Sorter100|10957_  = \new_Sorter100|10857_  & \new_Sorter100|10858_ ;
  assign \new_Sorter100|10958_  = \new_Sorter100|10857_  | \new_Sorter100|10858_ ;
  assign \new_Sorter100|10959_  = \new_Sorter100|10859_  & \new_Sorter100|10860_ ;
  assign \new_Sorter100|10960_  = \new_Sorter100|10859_  | \new_Sorter100|10860_ ;
  assign \new_Sorter100|10961_  = \new_Sorter100|10861_  & \new_Sorter100|10862_ ;
  assign \new_Sorter100|10962_  = \new_Sorter100|10861_  | \new_Sorter100|10862_ ;
  assign \new_Sorter100|10963_  = \new_Sorter100|10863_  & \new_Sorter100|10864_ ;
  assign \new_Sorter100|10964_  = \new_Sorter100|10863_  | \new_Sorter100|10864_ ;
  assign \new_Sorter100|10965_  = \new_Sorter100|10865_  & \new_Sorter100|10866_ ;
  assign \new_Sorter100|10966_  = \new_Sorter100|10865_  | \new_Sorter100|10866_ ;
  assign \new_Sorter100|10967_  = \new_Sorter100|10867_  & \new_Sorter100|10868_ ;
  assign \new_Sorter100|10968_  = \new_Sorter100|10867_  | \new_Sorter100|10868_ ;
  assign \new_Sorter100|10969_  = \new_Sorter100|10869_  & \new_Sorter100|10870_ ;
  assign \new_Sorter100|10970_  = \new_Sorter100|10869_  | \new_Sorter100|10870_ ;
  assign \new_Sorter100|10971_  = \new_Sorter100|10871_  & \new_Sorter100|10872_ ;
  assign \new_Sorter100|10972_  = \new_Sorter100|10871_  | \new_Sorter100|10872_ ;
  assign \new_Sorter100|10973_  = \new_Sorter100|10873_  & \new_Sorter100|10874_ ;
  assign \new_Sorter100|10974_  = \new_Sorter100|10873_  | \new_Sorter100|10874_ ;
  assign \new_Sorter100|10975_  = \new_Sorter100|10875_  & \new_Sorter100|10876_ ;
  assign \new_Sorter100|10976_  = \new_Sorter100|10875_  | \new_Sorter100|10876_ ;
  assign \new_Sorter100|10977_  = \new_Sorter100|10877_  & \new_Sorter100|10878_ ;
  assign \new_Sorter100|10978_  = \new_Sorter100|10877_  | \new_Sorter100|10878_ ;
  assign \new_Sorter100|10979_  = \new_Sorter100|10879_  & \new_Sorter100|10880_ ;
  assign \new_Sorter100|10980_  = \new_Sorter100|10879_  | \new_Sorter100|10880_ ;
  assign \new_Sorter100|10981_  = \new_Sorter100|10881_  & \new_Sorter100|10882_ ;
  assign \new_Sorter100|10982_  = \new_Sorter100|10881_  | \new_Sorter100|10882_ ;
  assign \new_Sorter100|10983_  = \new_Sorter100|10883_  & \new_Sorter100|10884_ ;
  assign \new_Sorter100|10984_  = \new_Sorter100|10883_  | \new_Sorter100|10884_ ;
  assign \new_Sorter100|10985_  = \new_Sorter100|10885_  & \new_Sorter100|10886_ ;
  assign \new_Sorter100|10986_  = \new_Sorter100|10885_  | \new_Sorter100|10886_ ;
  assign \new_Sorter100|10987_  = \new_Sorter100|10887_  & \new_Sorter100|10888_ ;
  assign \new_Sorter100|10988_  = \new_Sorter100|10887_  | \new_Sorter100|10888_ ;
  assign \new_Sorter100|10989_  = \new_Sorter100|10889_  & \new_Sorter100|10890_ ;
  assign \new_Sorter100|10990_  = \new_Sorter100|10889_  | \new_Sorter100|10890_ ;
  assign \new_Sorter100|10991_  = \new_Sorter100|10891_  & \new_Sorter100|10892_ ;
  assign \new_Sorter100|10992_  = \new_Sorter100|10891_  | \new_Sorter100|10892_ ;
  assign \new_Sorter100|10993_  = \new_Sorter100|10893_  & \new_Sorter100|10894_ ;
  assign \new_Sorter100|10994_  = \new_Sorter100|10893_  | \new_Sorter100|10894_ ;
  assign \new_Sorter100|10995_  = \new_Sorter100|10895_  & \new_Sorter100|10896_ ;
  assign \new_Sorter100|10996_  = \new_Sorter100|10895_  | \new_Sorter100|10896_ ;
  assign \new_Sorter100|10997_  = \new_Sorter100|10897_  & \new_Sorter100|10898_ ;
  assign \new_Sorter100|10998_  = \new_Sorter100|10897_  | \new_Sorter100|10898_ ;
  assign \new_Sorter100|11000_  = \new_Sorter100|10900_  & \new_Sorter100|10901_ ;
  assign \new_Sorter100|11001_  = \new_Sorter100|10900_  | \new_Sorter100|10901_ ;
  assign \new_Sorter100|11002_  = \new_Sorter100|10902_  & \new_Sorter100|10903_ ;
  assign \new_Sorter100|11003_  = \new_Sorter100|10902_  | \new_Sorter100|10903_ ;
  assign \new_Sorter100|11004_  = \new_Sorter100|10904_  & \new_Sorter100|10905_ ;
  assign \new_Sorter100|11005_  = \new_Sorter100|10904_  | \new_Sorter100|10905_ ;
  assign \new_Sorter100|11006_  = \new_Sorter100|10906_  & \new_Sorter100|10907_ ;
  assign \new_Sorter100|11007_  = \new_Sorter100|10906_  | \new_Sorter100|10907_ ;
  assign \new_Sorter100|11008_  = \new_Sorter100|10908_  & \new_Sorter100|10909_ ;
  assign \new_Sorter100|11009_  = \new_Sorter100|10908_  | \new_Sorter100|10909_ ;
  assign \new_Sorter100|11010_  = \new_Sorter100|10910_  & \new_Sorter100|10911_ ;
  assign \new_Sorter100|11011_  = \new_Sorter100|10910_  | \new_Sorter100|10911_ ;
  assign \new_Sorter100|11012_  = \new_Sorter100|10912_  & \new_Sorter100|10913_ ;
  assign \new_Sorter100|11013_  = \new_Sorter100|10912_  | \new_Sorter100|10913_ ;
  assign \new_Sorter100|11014_  = \new_Sorter100|10914_  & \new_Sorter100|10915_ ;
  assign \new_Sorter100|11015_  = \new_Sorter100|10914_  | \new_Sorter100|10915_ ;
  assign \new_Sorter100|11016_  = \new_Sorter100|10916_  & \new_Sorter100|10917_ ;
  assign \new_Sorter100|11017_  = \new_Sorter100|10916_  | \new_Sorter100|10917_ ;
  assign \new_Sorter100|11018_  = \new_Sorter100|10918_  & \new_Sorter100|10919_ ;
  assign \new_Sorter100|11019_  = \new_Sorter100|10918_  | \new_Sorter100|10919_ ;
  assign \new_Sorter100|11020_  = \new_Sorter100|10920_  & \new_Sorter100|10921_ ;
  assign \new_Sorter100|11021_  = \new_Sorter100|10920_  | \new_Sorter100|10921_ ;
  assign \new_Sorter100|11022_  = \new_Sorter100|10922_  & \new_Sorter100|10923_ ;
  assign \new_Sorter100|11023_  = \new_Sorter100|10922_  | \new_Sorter100|10923_ ;
  assign \new_Sorter100|11024_  = \new_Sorter100|10924_  & \new_Sorter100|10925_ ;
  assign \new_Sorter100|11025_  = \new_Sorter100|10924_  | \new_Sorter100|10925_ ;
  assign \new_Sorter100|11026_  = \new_Sorter100|10926_  & \new_Sorter100|10927_ ;
  assign \new_Sorter100|11027_  = \new_Sorter100|10926_  | \new_Sorter100|10927_ ;
  assign \new_Sorter100|11028_  = \new_Sorter100|10928_  & \new_Sorter100|10929_ ;
  assign \new_Sorter100|11029_  = \new_Sorter100|10928_  | \new_Sorter100|10929_ ;
  assign \new_Sorter100|11030_  = \new_Sorter100|10930_  & \new_Sorter100|10931_ ;
  assign \new_Sorter100|11031_  = \new_Sorter100|10930_  | \new_Sorter100|10931_ ;
  assign \new_Sorter100|11032_  = \new_Sorter100|10932_  & \new_Sorter100|10933_ ;
  assign \new_Sorter100|11033_  = \new_Sorter100|10932_  | \new_Sorter100|10933_ ;
  assign \new_Sorter100|11034_  = \new_Sorter100|10934_  & \new_Sorter100|10935_ ;
  assign \new_Sorter100|11035_  = \new_Sorter100|10934_  | \new_Sorter100|10935_ ;
  assign \new_Sorter100|11036_  = \new_Sorter100|10936_  & \new_Sorter100|10937_ ;
  assign \new_Sorter100|11037_  = \new_Sorter100|10936_  | \new_Sorter100|10937_ ;
  assign \new_Sorter100|11038_  = \new_Sorter100|10938_  & \new_Sorter100|10939_ ;
  assign \new_Sorter100|11039_  = \new_Sorter100|10938_  | \new_Sorter100|10939_ ;
  assign \new_Sorter100|11040_  = \new_Sorter100|10940_  & \new_Sorter100|10941_ ;
  assign \new_Sorter100|11041_  = \new_Sorter100|10940_  | \new_Sorter100|10941_ ;
  assign \new_Sorter100|11042_  = \new_Sorter100|10942_  & \new_Sorter100|10943_ ;
  assign \new_Sorter100|11043_  = \new_Sorter100|10942_  | \new_Sorter100|10943_ ;
  assign \new_Sorter100|11044_  = \new_Sorter100|10944_  & \new_Sorter100|10945_ ;
  assign \new_Sorter100|11045_  = \new_Sorter100|10944_  | \new_Sorter100|10945_ ;
  assign \new_Sorter100|11046_  = \new_Sorter100|10946_  & \new_Sorter100|10947_ ;
  assign \new_Sorter100|11047_  = \new_Sorter100|10946_  | \new_Sorter100|10947_ ;
  assign \new_Sorter100|11048_  = \new_Sorter100|10948_  & \new_Sorter100|10949_ ;
  assign \new_Sorter100|11049_  = \new_Sorter100|10948_  | \new_Sorter100|10949_ ;
  assign \new_Sorter100|11050_  = \new_Sorter100|10950_  & \new_Sorter100|10951_ ;
  assign \new_Sorter100|11051_  = \new_Sorter100|10950_  | \new_Sorter100|10951_ ;
  assign \new_Sorter100|11052_  = \new_Sorter100|10952_  & \new_Sorter100|10953_ ;
  assign \new_Sorter100|11053_  = \new_Sorter100|10952_  | \new_Sorter100|10953_ ;
  assign \new_Sorter100|11054_  = \new_Sorter100|10954_  & \new_Sorter100|10955_ ;
  assign \new_Sorter100|11055_  = \new_Sorter100|10954_  | \new_Sorter100|10955_ ;
  assign \new_Sorter100|11056_  = \new_Sorter100|10956_  & \new_Sorter100|10957_ ;
  assign \new_Sorter100|11057_  = \new_Sorter100|10956_  | \new_Sorter100|10957_ ;
  assign \new_Sorter100|11058_  = \new_Sorter100|10958_  & \new_Sorter100|10959_ ;
  assign \new_Sorter100|11059_  = \new_Sorter100|10958_  | \new_Sorter100|10959_ ;
  assign \new_Sorter100|11060_  = \new_Sorter100|10960_  & \new_Sorter100|10961_ ;
  assign \new_Sorter100|11061_  = \new_Sorter100|10960_  | \new_Sorter100|10961_ ;
  assign \new_Sorter100|11062_  = \new_Sorter100|10962_  & \new_Sorter100|10963_ ;
  assign \new_Sorter100|11063_  = \new_Sorter100|10962_  | \new_Sorter100|10963_ ;
  assign \new_Sorter100|11064_  = \new_Sorter100|10964_  & \new_Sorter100|10965_ ;
  assign \new_Sorter100|11065_  = \new_Sorter100|10964_  | \new_Sorter100|10965_ ;
  assign \new_Sorter100|11066_  = \new_Sorter100|10966_  & \new_Sorter100|10967_ ;
  assign \new_Sorter100|11067_  = \new_Sorter100|10966_  | \new_Sorter100|10967_ ;
  assign \new_Sorter100|11068_  = \new_Sorter100|10968_  & \new_Sorter100|10969_ ;
  assign \new_Sorter100|11069_  = \new_Sorter100|10968_  | \new_Sorter100|10969_ ;
  assign \new_Sorter100|11070_  = \new_Sorter100|10970_  & \new_Sorter100|10971_ ;
  assign \new_Sorter100|11071_  = \new_Sorter100|10970_  | \new_Sorter100|10971_ ;
  assign \new_Sorter100|11072_  = \new_Sorter100|10972_  & \new_Sorter100|10973_ ;
  assign \new_Sorter100|11073_  = \new_Sorter100|10972_  | \new_Sorter100|10973_ ;
  assign \new_Sorter100|11074_  = \new_Sorter100|10974_  & \new_Sorter100|10975_ ;
  assign \new_Sorter100|11075_  = \new_Sorter100|10974_  | \new_Sorter100|10975_ ;
  assign \new_Sorter100|11076_  = \new_Sorter100|10976_  & \new_Sorter100|10977_ ;
  assign \new_Sorter100|11077_  = \new_Sorter100|10976_  | \new_Sorter100|10977_ ;
  assign \new_Sorter100|11078_  = \new_Sorter100|10978_  & \new_Sorter100|10979_ ;
  assign \new_Sorter100|11079_  = \new_Sorter100|10978_  | \new_Sorter100|10979_ ;
  assign \new_Sorter100|11080_  = \new_Sorter100|10980_  & \new_Sorter100|10981_ ;
  assign \new_Sorter100|11081_  = \new_Sorter100|10980_  | \new_Sorter100|10981_ ;
  assign \new_Sorter100|11082_  = \new_Sorter100|10982_  & \new_Sorter100|10983_ ;
  assign \new_Sorter100|11083_  = \new_Sorter100|10982_  | \new_Sorter100|10983_ ;
  assign \new_Sorter100|11084_  = \new_Sorter100|10984_  & \new_Sorter100|10985_ ;
  assign \new_Sorter100|11085_  = \new_Sorter100|10984_  | \new_Sorter100|10985_ ;
  assign \new_Sorter100|11086_  = \new_Sorter100|10986_  & \new_Sorter100|10987_ ;
  assign \new_Sorter100|11087_  = \new_Sorter100|10986_  | \new_Sorter100|10987_ ;
  assign \new_Sorter100|11088_  = \new_Sorter100|10988_  & \new_Sorter100|10989_ ;
  assign \new_Sorter100|11089_  = \new_Sorter100|10988_  | \new_Sorter100|10989_ ;
  assign \new_Sorter100|11090_  = \new_Sorter100|10990_  & \new_Sorter100|10991_ ;
  assign \new_Sorter100|11091_  = \new_Sorter100|10990_  | \new_Sorter100|10991_ ;
  assign \new_Sorter100|11092_  = \new_Sorter100|10992_  & \new_Sorter100|10993_ ;
  assign \new_Sorter100|11093_  = \new_Sorter100|10992_  | \new_Sorter100|10993_ ;
  assign \new_Sorter100|11094_  = \new_Sorter100|10994_  & \new_Sorter100|10995_ ;
  assign \new_Sorter100|11095_  = \new_Sorter100|10994_  | \new_Sorter100|10995_ ;
  assign \new_Sorter100|11096_  = \new_Sorter100|10996_  & \new_Sorter100|10997_ ;
  assign \new_Sorter100|11097_  = \new_Sorter100|10996_  | \new_Sorter100|10997_ ;
  assign \new_Sorter100|11098_  = \new_Sorter100|10998_  & \new_Sorter100|10999_ ;
  assign \new_Sorter100|11099_  = \new_Sorter100|10998_  | \new_Sorter100|10999_ ;
  assign \new_Sorter100|11100_  = \new_Sorter100|11000_ ;
  assign \new_Sorter100|11199_  = \new_Sorter100|11099_ ;
  assign \new_Sorter100|11101_  = \new_Sorter100|11001_  & \new_Sorter100|11002_ ;
  assign \new_Sorter100|11102_  = \new_Sorter100|11001_  | \new_Sorter100|11002_ ;
  assign \new_Sorter100|11103_  = \new_Sorter100|11003_  & \new_Sorter100|11004_ ;
  assign \new_Sorter100|11104_  = \new_Sorter100|11003_  | \new_Sorter100|11004_ ;
  assign \new_Sorter100|11105_  = \new_Sorter100|11005_  & \new_Sorter100|11006_ ;
  assign \new_Sorter100|11106_  = \new_Sorter100|11005_  | \new_Sorter100|11006_ ;
  assign \new_Sorter100|11107_  = \new_Sorter100|11007_  & \new_Sorter100|11008_ ;
  assign \new_Sorter100|11108_  = \new_Sorter100|11007_  | \new_Sorter100|11008_ ;
  assign \new_Sorter100|11109_  = \new_Sorter100|11009_  & \new_Sorter100|11010_ ;
  assign \new_Sorter100|11110_  = \new_Sorter100|11009_  | \new_Sorter100|11010_ ;
  assign \new_Sorter100|11111_  = \new_Sorter100|11011_  & \new_Sorter100|11012_ ;
  assign \new_Sorter100|11112_  = \new_Sorter100|11011_  | \new_Sorter100|11012_ ;
  assign \new_Sorter100|11113_  = \new_Sorter100|11013_  & \new_Sorter100|11014_ ;
  assign \new_Sorter100|11114_  = \new_Sorter100|11013_  | \new_Sorter100|11014_ ;
  assign \new_Sorter100|11115_  = \new_Sorter100|11015_  & \new_Sorter100|11016_ ;
  assign \new_Sorter100|11116_  = \new_Sorter100|11015_  | \new_Sorter100|11016_ ;
  assign \new_Sorter100|11117_  = \new_Sorter100|11017_  & \new_Sorter100|11018_ ;
  assign \new_Sorter100|11118_  = \new_Sorter100|11017_  | \new_Sorter100|11018_ ;
  assign \new_Sorter100|11119_  = \new_Sorter100|11019_  & \new_Sorter100|11020_ ;
  assign \new_Sorter100|11120_  = \new_Sorter100|11019_  | \new_Sorter100|11020_ ;
  assign \new_Sorter100|11121_  = \new_Sorter100|11021_  & \new_Sorter100|11022_ ;
  assign \new_Sorter100|11122_  = \new_Sorter100|11021_  | \new_Sorter100|11022_ ;
  assign \new_Sorter100|11123_  = \new_Sorter100|11023_  & \new_Sorter100|11024_ ;
  assign \new_Sorter100|11124_  = \new_Sorter100|11023_  | \new_Sorter100|11024_ ;
  assign \new_Sorter100|11125_  = \new_Sorter100|11025_  & \new_Sorter100|11026_ ;
  assign \new_Sorter100|11126_  = \new_Sorter100|11025_  | \new_Sorter100|11026_ ;
  assign \new_Sorter100|11127_  = \new_Sorter100|11027_  & \new_Sorter100|11028_ ;
  assign \new_Sorter100|11128_  = \new_Sorter100|11027_  | \new_Sorter100|11028_ ;
  assign \new_Sorter100|11129_  = \new_Sorter100|11029_  & \new_Sorter100|11030_ ;
  assign \new_Sorter100|11130_  = \new_Sorter100|11029_  | \new_Sorter100|11030_ ;
  assign \new_Sorter100|11131_  = \new_Sorter100|11031_  & \new_Sorter100|11032_ ;
  assign \new_Sorter100|11132_  = \new_Sorter100|11031_  | \new_Sorter100|11032_ ;
  assign \new_Sorter100|11133_  = \new_Sorter100|11033_  & \new_Sorter100|11034_ ;
  assign \new_Sorter100|11134_  = \new_Sorter100|11033_  | \new_Sorter100|11034_ ;
  assign \new_Sorter100|11135_  = \new_Sorter100|11035_  & \new_Sorter100|11036_ ;
  assign \new_Sorter100|11136_  = \new_Sorter100|11035_  | \new_Sorter100|11036_ ;
  assign \new_Sorter100|11137_  = \new_Sorter100|11037_  & \new_Sorter100|11038_ ;
  assign \new_Sorter100|11138_  = \new_Sorter100|11037_  | \new_Sorter100|11038_ ;
  assign \new_Sorter100|11139_  = \new_Sorter100|11039_  & \new_Sorter100|11040_ ;
  assign \new_Sorter100|11140_  = \new_Sorter100|11039_  | \new_Sorter100|11040_ ;
  assign \new_Sorter100|11141_  = \new_Sorter100|11041_  & \new_Sorter100|11042_ ;
  assign \new_Sorter100|11142_  = \new_Sorter100|11041_  | \new_Sorter100|11042_ ;
  assign \new_Sorter100|11143_  = \new_Sorter100|11043_  & \new_Sorter100|11044_ ;
  assign \new_Sorter100|11144_  = \new_Sorter100|11043_  | \new_Sorter100|11044_ ;
  assign \new_Sorter100|11145_  = \new_Sorter100|11045_  & \new_Sorter100|11046_ ;
  assign \new_Sorter100|11146_  = \new_Sorter100|11045_  | \new_Sorter100|11046_ ;
  assign \new_Sorter100|11147_  = \new_Sorter100|11047_  & \new_Sorter100|11048_ ;
  assign \new_Sorter100|11148_  = \new_Sorter100|11047_  | \new_Sorter100|11048_ ;
  assign \new_Sorter100|11149_  = \new_Sorter100|11049_  & \new_Sorter100|11050_ ;
  assign \new_Sorter100|11150_  = \new_Sorter100|11049_  | \new_Sorter100|11050_ ;
  assign \new_Sorter100|11151_  = \new_Sorter100|11051_  & \new_Sorter100|11052_ ;
  assign \new_Sorter100|11152_  = \new_Sorter100|11051_  | \new_Sorter100|11052_ ;
  assign \new_Sorter100|11153_  = \new_Sorter100|11053_  & \new_Sorter100|11054_ ;
  assign \new_Sorter100|11154_  = \new_Sorter100|11053_  | \new_Sorter100|11054_ ;
  assign \new_Sorter100|11155_  = \new_Sorter100|11055_  & \new_Sorter100|11056_ ;
  assign \new_Sorter100|11156_  = \new_Sorter100|11055_  | \new_Sorter100|11056_ ;
  assign \new_Sorter100|11157_  = \new_Sorter100|11057_  & \new_Sorter100|11058_ ;
  assign \new_Sorter100|11158_  = \new_Sorter100|11057_  | \new_Sorter100|11058_ ;
  assign \new_Sorter100|11159_  = \new_Sorter100|11059_  & \new_Sorter100|11060_ ;
  assign \new_Sorter100|11160_  = \new_Sorter100|11059_  | \new_Sorter100|11060_ ;
  assign \new_Sorter100|11161_  = \new_Sorter100|11061_  & \new_Sorter100|11062_ ;
  assign \new_Sorter100|11162_  = \new_Sorter100|11061_  | \new_Sorter100|11062_ ;
  assign \new_Sorter100|11163_  = \new_Sorter100|11063_  & \new_Sorter100|11064_ ;
  assign \new_Sorter100|11164_  = \new_Sorter100|11063_  | \new_Sorter100|11064_ ;
  assign \new_Sorter100|11165_  = \new_Sorter100|11065_  & \new_Sorter100|11066_ ;
  assign \new_Sorter100|11166_  = \new_Sorter100|11065_  | \new_Sorter100|11066_ ;
  assign \new_Sorter100|11167_  = \new_Sorter100|11067_  & \new_Sorter100|11068_ ;
  assign \new_Sorter100|11168_  = \new_Sorter100|11067_  | \new_Sorter100|11068_ ;
  assign \new_Sorter100|11169_  = \new_Sorter100|11069_  & \new_Sorter100|11070_ ;
  assign \new_Sorter100|11170_  = \new_Sorter100|11069_  | \new_Sorter100|11070_ ;
  assign \new_Sorter100|11171_  = \new_Sorter100|11071_  & \new_Sorter100|11072_ ;
  assign \new_Sorter100|11172_  = \new_Sorter100|11071_  | \new_Sorter100|11072_ ;
  assign \new_Sorter100|11173_  = \new_Sorter100|11073_  & \new_Sorter100|11074_ ;
  assign \new_Sorter100|11174_  = \new_Sorter100|11073_  | \new_Sorter100|11074_ ;
  assign \new_Sorter100|11175_  = \new_Sorter100|11075_  & \new_Sorter100|11076_ ;
  assign \new_Sorter100|11176_  = \new_Sorter100|11075_  | \new_Sorter100|11076_ ;
  assign \new_Sorter100|11177_  = \new_Sorter100|11077_  & \new_Sorter100|11078_ ;
  assign \new_Sorter100|11178_  = \new_Sorter100|11077_  | \new_Sorter100|11078_ ;
  assign \new_Sorter100|11179_  = \new_Sorter100|11079_  & \new_Sorter100|11080_ ;
  assign \new_Sorter100|11180_  = \new_Sorter100|11079_  | \new_Sorter100|11080_ ;
  assign \new_Sorter100|11181_  = \new_Sorter100|11081_  & \new_Sorter100|11082_ ;
  assign \new_Sorter100|11182_  = \new_Sorter100|11081_  | \new_Sorter100|11082_ ;
  assign \new_Sorter100|11183_  = \new_Sorter100|11083_  & \new_Sorter100|11084_ ;
  assign \new_Sorter100|11184_  = \new_Sorter100|11083_  | \new_Sorter100|11084_ ;
  assign \new_Sorter100|11185_  = \new_Sorter100|11085_  & \new_Sorter100|11086_ ;
  assign \new_Sorter100|11186_  = \new_Sorter100|11085_  | \new_Sorter100|11086_ ;
  assign \new_Sorter100|11187_  = \new_Sorter100|11087_  & \new_Sorter100|11088_ ;
  assign \new_Sorter100|11188_  = \new_Sorter100|11087_  | \new_Sorter100|11088_ ;
  assign \new_Sorter100|11189_  = \new_Sorter100|11089_  & \new_Sorter100|11090_ ;
  assign \new_Sorter100|11190_  = \new_Sorter100|11089_  | \new_Sorter100|11090_ ;
  assign \new_Sorter100|11191_  = \new_Sorter100|11091_  & \new_Sorter100|11092_ ;
  assign \new_Sorter100|11192_  = \new_Sorter100|11091_  | \new_Sorter100|11092_ ;
  assign \new_Sorter100|11193_  = \new_Sorter100|11093_  & \new_Sorter100|11094_ ;
  assign \new_Sorter100|11194_  = \new_Sorter100|11093_  | \new_Sorter100|11094_ ;
  assign \new_Sorter100|11195_  = \new_Sorter100|11095_  & \new_Sorter100|11096_ ;
  assign \new_Sorter100|11196_  = \new_Sorter100|11095_  | \new_Sorter100|11096_ ;
  assign \new_Sorter100|11197_  = \new_Sorter100|11097_  & \new_Sorter100|11098_ ;
  assign \new_Sorter100|11198_  = \new_Sorter100|11097_  | \new_Sorter100|11098_ ;
  assign \new_Sorter100|11200_  = \new_Sorter100|11100_  & \new_Sorter100|11101_ ;
  assign \new_Sorter100|11201_  = \new_Sorter100|11100_  | \new_Sorter100|11101_ ;
  assign \new_Sorter100|11202_  = \new_Sorter100|11102_  & \new_Sorter100|11103_ ;
  assign \new_Sorter100|11203_  = \new_Sorter100|11102_  | \new_Sorter100|11103_ ;
  assign \new_Sorter100|11204_  = \new_Sorter100|11104_  & \new_Sorter100|11105_ ;
  assign \new_Sorter100|11205_  = \new_Sorter100|11104_  | \new_Sorter100|11105_ ;
  assign \new_Sorter100|11206_  = \new_Sorter100|11106_  & \new_Sorter100|11107_ ;
  assign \new_Sorter100|11207_  = \new_Sorter100|11106_  | \new_Sorter100|11107_ ;
  assign \new_Sorter100|11208_  = \new_Sorter100|11108_  & \new_Sorter100|11109_ ;
  assign \new_Sorter100|11209_  = \new_Sorter100|11108_  | \new_Sorter100|11109_ ;
  assign \new_Sorter100|11210_  = \new_Sorter100|11110_  & \new_Sorter100|11111_ ;
  assign \new_Sorter100|11211_  = \new_Sorter100|11110_  | \new_Sorter100|11111_ ;
  assign \new_Sorter100|11212_  = \new_Sorter100|11112_  & \new_Sorter100|11113_ ;
  assign \new_Sorter100|11213_  = \new_Sorter100|11112_  | \new_Sorter100|11113_ ;
  assign \new_Sorter100|11214_  = \new_Sorter100|11114_  & \new_Sorter100|11115_ ;
  assign \new_Sorter100|11215_  = \new_Sorter100|11114_  | \new_Sorter100|11115_ ;
  assign \new_Sorter100|11216_  = \new_Sorter100|11116_  & \new_Sorter100|11117_ ;
  assign \new_Sorter100|11217_  = \new_Sorter100|11116_  | \new_Sorter100|11117_ ;
  assign \new_Sorter100|11218_  = \new_Sorter100|11118_  & \new_Sorter100|11119_ ;
  assign \new_Sorter100|11219_  = \new_Sorter100|11118_  | \new_Sorter100|11119_ ;
  assign \new_Sorter100|11220_  = \new_Sorter100|11120_  & \new_Sorter100|11121_ ;
  assign \new_Sorter100|11221_  = \new_Sorter100|11120_  | \new_Sorter100|11121_ ;
  assign \new_Sorter100|11222_  = \new_Sorter100|11122_  & \new_Sorter100|11123_ ;
  assign \new_Sorter100|11223_  = \new_Sorter100|11122_  | \new_Sorter100|11123_ ;
  assign \new_Sorter100|11224_  = \new_Sorter100|11124_  & \new_Sorter100|11125_ ;
  assign \new_Sorter100|11225_  = \new_Sorter100|11124_  | \new_Sorter100|11125_ ;
  assign \new_Sorter100|11226_  = \new_Sorter100|11126_  & \new_Sorter100|11127_ ;
  assign \new_Sorter100|11227_  = \new_Sorter100|11126_  | \new_Sorter100|11127_ ;
  assign \new_Sorter100|11228_  = \new_Sorter100|11128_  & \new_Sorter100|11129_ ;
  assign \new_Sorter100|11229_  = \new_Sorter100|11128_  | \new_Sorter100|11129_ ;
  assign \new_Sorter100|11230_  = \new_Sorter100|11130_  & \new_Sorter100|11131_ ;
  assign \new_Sorter100|11231_  = \new_Sorter100|11130_  | \new_Sorter100|11131_ ;
  assign \new_Sorter100|11232_  = \new_Sorter100|11132_  & \new_Sorter100|11133_ ;
  assign \new_Sorter100|11233_  = \new_Sorter100|11132_  | \new_Sorter100|11133_ ;
  assign \new_Sorter100|11234_  = \new_Sorter100|11134_  & \new_Sorter100|11135_ ;
  assign \new_Sorter100|11235_  = \new_Sorter100|11134_  | \new_Sorter100|11135_ ;
  assign \new_Sorter100|11236_  = \new_Sorter100|11136_  & \new_Sorter100|11137_ ;
  assign \new_Sorter100|11237_  = \new_Sorter100|11136_  | \new_Sorter100|11137_ ;
  assign \new_Sorter100|11238_  = \new_Sorter100|11138_  & \new_Sorter100|11139_ ;
  assign \new_Sorter100|11239_  = \new_Sorter100|11138_  | \new_Sorter100|11139_ ;
  assign \new_Sorter100|11240_  = \new_Sorter100|11140_  & \new_Sorter100|11141_ ;
  assign \new_Sorter100|11241_  = \new_Sorter100|11140_  | \new_Sorter100|11141_ ;
  assign \new_Sorter100|11242_  = \new_Sorter100|11142_  & \new_Sorter100|11143_ ;
  assign \new_Sorter100|11243_  = \new_Sorter100|11142_  | \new_Sorter100|11143_ ;
  assign \new_Sorter100|11244_  = \new_Sorter100|11144_  & \new_Sorter100|11145_ ;
  assign \new_Sorter100|11245_  = \new_Sorter100|11144_  | \new_Sorter100|11145_ ;
  assign \new_Sorter100|11246_  = \new_Sorter100|11146_  & \new_Sorter100|11147_ ;
  assign \new_Sorter100|11247_  = \new_Sorter100|11146_  | \new_Sorter100|11147_ ;
  assign \new_Sorter100|11248_  = \new_Sorter100|11148_  & \new_Sorter100|11149_ ;
  assign \new_Sorter100|11249_  = \new_Sorter100|11148_  | \new_Sorter100|11149_ ;
  assign \new_Sorter100|11250_  = \new_Sorter100|11150_  & \new_Sorter100|11151_ ;
  assign \new_Sorter100|11251_  = \new_Sorter100|11150_  | \new_Sorter100|11151_ ;
  assign \new_Sorter100|11252_  = \new_Sorter100|11152_  & \new_Sorter100|11153_ ;
  assign \new_Sorter100|11253_  = \new_Sorter100|11152_  | \new_Sorter100|11153_ ;
  assign \new_Sorter100|11254_  = \new_Sorter100|11154_  & \new_Sorter100|11155_ ;
  assign \new_Sorter100|11255_  = \new_Sorter100|11154_  | \new_Sorter100|11155_ ;
  assign \new_Sorter100|11256_  = \new_Sorter100|11156_  & \new_Sorter100|11157_ ;
  assign \new_Sorter100|11257_  = \new_Sorter100|11156_  | \new_Sorter100|11157_ ;
  assign \new_Sorter100|11258_  = \new_Sorter100|11158_  & \new_Sorter100|11159_ ;
  assign \new_Sorter100|11259_  = \new_Sorter100|11158_  | \new_Sorter100|11159_ ;
  assign \new_Sorter100|11260_  = \new_Sorter100|11160_  & \new_Sorter100|11161_ ;
  assign \new_Sorter100|11261_  = \new_Sorter100|11160_  | \new_Sorter100|11161_ ;
  assign \new_Sorter100|11262_  = \new_Sorter100|11162_  & \new_Sorter100|11163_ ;
  assign \new_Sorter100|11263_  = \new_Sorter100|11162_  | \new_Sorter100|11163_ ;
  assign \new_Sorter100|11264_  = \new_Sorter100|11164_  & \new_Sorter100|11165_ ;
  assign \new_Sorter100|11265_  = \new_Sorter100|11164_  | \new_Sorter100|11165_ ;
  assign \new_Sorter100|11266_  = \new_Sorter100|11166_  & \new_Sorter100|11167_ ;
  assign \new_Sorter100|11267_  = \new_Sorter100|11166_  | \new_Sorter100|11167_ ;
  assign \new_Sorter100|11268_  = \new_Sorter100|11168_  & \new_Sorter100|11169_ ;
  assign \new_Sorter100|11269_  = \new_Sorter100|11168_  | \new_Sorter100|11169_ ;
  assign \new_Sorter100|11270_  = \new_Sorter100|11170_  & \new_Sorter100|11171_ ;
  assign \new_Sorter100|11271_  = \new_Sorter100|11170_  | \new_Sorter100|11171_ ;
  assign \new_Sorter100|11272_  = \new_Sorter100|11172_  & \new_Sorter100|11173_ ;
  assign \new_Sorter100|11273_  = \new_Sorter100|11172_  | \new_Sorter100|11173_ ;
  assign \new_Sorter100|11274_  = \new_Sorter100|11174_  & \new_Sorter100|11175_ ;
  assign \new_Sorter100|11275_  = \new_Sorter100|11174_  | \new_Sorter100|11175_ ;
  assign \new_Sorter100|11276_  = \new_Sorter100|11176_  & \new_Sorter100|11177_ ;
  assign \new_Sorter100|11277_  = \new_Sorter100|11176_  | \new_Sorter100|11177_ ;
  assign \new_Sorter100|11278_  = \new_Sorter100|11178_  & \new_Sorter100|11179_ ;
  assign \new_Sorter100|11279_  = \new_Sorter100|11178_  | \new_Sorter100|11179_ ;
  assign \new_Sorter100|11280_  = \new_Sorter100|11180_  & \new_Sorter100|11181_ ;
  assign \new_Sorter100|11281_  = \new_Sorter100|11180_  | \new_Sorter100|11181_ ;
  assign \new_Sorter100|11282_  = \new_Sorter100|11182_  & \new_Sorter100|11183_ ;
  assign \new_Sorter100|11283_  = \new_Sorter100|11182_  | \new_Sorter100|11183_ ;
  assign \new_Sorter100|11284_  = \new_Sorter100|11184_  & \new_Sorter100|11185_ ;
  assign \new_Sorter100|11285_  = \new_Sorter100|11184_  | \new_Sorter100|11185_ ;
  assign \new_Sorter100|11286_  = \new_Sorter100|11186_  & \new_Sorter100|11187_ ;
  assign \new_Sorter100|11287_  = \new_Sorter100|11186_  | \new_Sorter100|11187_ ;
  assign \new_Sorter100|11288_  = \new_Sorter100|11188_  & \new_Sorter100|11189_ ;
  assign \new_Sorter100|11289_  = \new_Sorter100|11188_  | \new_Sorter100|11189_ ;
  assign \new_Sorter100|11290_  = \new_Sorter100|11190_  & \new_Sorter100|11191_ ;
  assign \new_Sorter100|11291_  = \new_Sorter100|11190_  | \new_Sorter100|11191_ ;
  assign \new_Sorter100|11292_  = \new_Sorter100|11192_  & \new_Sorter100|11193_ ;
  assign \new_Sorter100|11293_  = \new_Sorter100|11192_  | \new_Sorter100|11193_ ;
  assign \new_Sorter100|11294_  = \new_Sorter100|11194_  & \new_Sorter100|11195_ ;
  assign \new_Sorter100|11295_  = \new_Sorter100|11194_  | \new_Sorter100|11195_ ;
  assign \new_Sorter100|11296_  = \new_Sorter100|11196_  & \new_Sorter100|11197_ ;
  assign \new_Sorter100|11297_  = \new_Sorter100|11196_  | \new_Sorter100|11197_ ;
  assign \new_Sorter100|11298_  = \new_Sorter100|11198_  & \new_Sorter100|11199_ ;
  assign \new_Sorter100|11299_  = \new_Sorter100|11198_  | \new_Sorter100|11199_ ;
  assign \new_Sorter100|11300_  = \new_Sorter100|11200_ ;
  assign \new_Sorter100|11399_  = \new_Sorter100|11299_ ;
  assign \new_Sorter100|11301_  = \new_Sorter100|11201_  & \new_Sorter100|11202_ ;
  assign \new_Sorter100|11302_  = \new_Sorter100|11201_  | \new_Sorter100|11202_ ;
  assign \new_Sorter100|11303_  = \new_Sorter100|11203_  & \new_Sorter100|11204_ ;
  assign \new_Sorter100|11304_  = \new_Sorter100|11203_  | \new_Sorter100|11204_ ;
  assign \new_Sorter100|11305_  = \new_Sorter100|11205_  & \new_Sorter100|11206_ ;
  assign \new_Sorter100|11306_  = \new_Sorter100|11205_  | \new_Sorter100|11206_ ;
  assign \new_Sorter100|11307_  = \new_Sorter100|11207_  & \new_Sorter100|11208_ ;
  assign \new_Sorter100|11308_  = \new_Sorter100|11207_  | \new_Sorter100|11208_ ;
  assign \new_Sorter100|11309_  = \new_Sorter100|11209_  & \new_Sorter100|11210_ ;
  assign \new_Sorter100|11310_  = \new_Sorter100|11209_  | \new_Sorter100|11210_ ;
  assign \new_Sorter100|11311_  = \new_Sorter100|11211_  & \new_Sorter100|11212_ ;
  assign \new_Sorter100|11312_  = \new_Sorter100|11211_  | \new_Sorter100|11212_ ;
  assign \new_Sorter100|11313_  = \new_Sorter100|11213_  & \new_Sorter100|11214_ ;
  assign \new_Sorter100|11314_  = \new_Sorter100|11213_  | \new_Sorter100|11214_ ;
  assign \new_Sorter100|11315_  = \new_Sorter100|11215_  & \new_Sorter100|11216_ ;
  assign \new_Sorter100|11316_  = \new_Sorter100|11215_  | \new_Sorter100|11216_ ;
  assign \new_Sorter100|11317_  = \new_Sorter100|11217_  & \new_Sorter100|11218_ ;
  assign \new_Sorter100|11318_  = \new_Sorter100|11217_  | \new_Sorter100|11218_ ;
  assign \new_Sorter100|11319_  = \new_Sorter100|11219_  & \new_Sorter100|11220_ ;
  assign \new_Sorter100|11320_  = \new_Sorter100|11219_  | \new_Sorter100|11220_ ;
  assign \new_Sorter100|11321_  = \new_Sorter100|11221_  & \new_Sorter100|11222_ ;
  assign \new_Sorter100|11322_  = \new_Sorter100|11221_  | \new_Sorter100|11222_ ;
  assign \new_Sorter100|11323_  = \new_Sorter100|11223_  & \new_Sorter100|11224_ ;
  assign \new_Sorter100|11324_  = \new_Sorter100|11223_  | \new_Sorter100|11224_ ;
  assign \new_Sorter100|11325_  = \new_Sorter100|11225_  & \new_Sorter100|11226_ ;
  assign \new_Sorter100|11326_  = \new_Sorter100|11225_  | \new_Sorter100|11226_ ;
  assign \new_Sorter100|11327_  = \new_Sorter100|11227_  & \new_Sorter100|11228_ ;
  assign \new_Sorter100|11328_  = \new_Sorter100|11227_  | \new_Sorter100|11228_ ;
  assign \new_Sorter100|11329_  = \new_Sorter100|11229_  & \new_Sorter100|11230_ ;
  assign \new_Sorter100|11330_  = \new_Sorter100|11229_  | \new_Sorter100|11230_ ;
  assign \new_Sorter100|11331_  = \new_Sorter100|11231_  & \new_Sorter100|11232_ ;
  assign \new_Sorter100|11332_  = \new_Sorter100|11231_  | \new_Sorter100|11232_ ;
  assign \new_Sorter100|11333_  = \new_Sorter100|11233_  & \new_Sorter100|11234_ ;
  assign \new_Sorter100|11334_  = \new_Sorter100|11233_  | \new_Sorter100|11234_ ;
  assign \new_Sorter100|11335_  = \new_Sorter100|11235_  & \new_Sorter100|11236_ ;
  assign \new_Sorter100|11336_  = \new_Sorter100|11235_  | \new_Sorter100|11236_ ;
  assign \new_Sorter100|11337_  = \new_Sorter100|11237_  & \new_Sorter100|11238_ ;
  assign \new_Sorter100|11338_  = \new_Sorter100|11237_  | \new_Sorter100|11238_ ;
  assign \new_Sorter100|11339_  = \new_Sorter100|11239_  & \new_Sorter100|11240_ ;
  assign \new_Sorter100|11340_  = \new_Sorter100|11239_  | \new_Sorter100|11240_ ;
  assign \new_Sorter100|11341_  = \new_Sorter100|11241_  & \new_Sorter100|11242_ ;
  assign \new_Sorter100|11342_  = \new_Sorter100|11241_  | \new_Sorter100|11242_ ;
  assign \new_Sorter100|11343_  = \new_Sorter100|11243_  & \new_Sorter100|11244_ ;
  assign \new_Sorter100|11344_  = \new_Sorter100|11243_  | \new_Sorter100|11244_ ;
  assign \new_Sorter100|11345_  = \new_Sorter100|11245_  & \new_Sorter100|11246_ ;
  assign \new_Sorter100|11346_  = \new_Sorter100|11245_  | \new_Sorter100|11246_ ;
  assign \new_Sorter100|11347_  = \new_Sorter100|11247_  & \new_Sorter100|11248_ ;
  assign \new_Sorter100|11348_  = \new_Sorter100|11247_  | \new_Sorter100|11248_ ;
  assign \new_Sorter100|11349_  = \new_Sorter100|11249_  & \new_Sorter100|11250_ ;
  assign \new_Sorter100|11350_  = \new_Sorter100|11249_  | \new_Sorter100|11250_ ;
  assign \new_Sorter100|11351_  = \new_Sorter100|11251_  & \new_Sorter100|11252_ ;
  assign \new_Sorter100|11352_  = \new_Sorter100|11251_  | \new_Sorter100|11252_ ;
  assign \new_Sorter100|11353_  = \new_Sorter100|11253_  & \new_Sorter100|11254_ ;
  assign \new_Sorter100|11354_  = \new_Sorter100|11253_  | \new_Sorter100|11254_ ;
  assign \new_Sorter100|11355_  = \new_Sorter100|11255_  & \new_Sorter100|11256_ ;
  assign \new_Sorter100|11356_  = \new_Sorter100|11255_  | \new_Sorter100|11256_ ;
  assign \new_Sorter100|11357_  = \new_Sorter100|11257_  & \new_Sorter100|11258_ ;
  assign \new_Sorter100|11358_  = \new_Sorter100|11257_  | \new_Sorter100|11258_ ;
  assign \new_Sorter100|11359_  = \new_Sorter100|11259_  & \new_Sorter100|11260_ ;
  assign \new_Sorter100|11360_  = \new_Sorter100|11259_  | \new_Sorter100|11260_ ;
  assign \new_Sorter100|11361_  = \new_Sorter100|11261_  & \new_Sorter100|11262_ ;
  assign \new_Sorter100|11362_  = \new_Sorter100|11261_  | \new_Sorter100|11262_ ;
  assign \new_Sorter100|11363_  = \new_Sorter100|11263_  & \new_Sorter100|11264_ ;
  assign \new_Sorter100|11364_  = \new_Sorter100|11263_  | \new_Sorter100|11264_ ;
  assign \new_Sorter100|11365_  = \new_Sorter100|11265_  & \new_Sorter100|11266_ ;
  assign \new_Sorter100|11366_  = \new_Sorter100|11265_  | \new_Sorter100|11266_ ;
  assign \new_Sorter100|11367_  = \new_Sorter100|11267_  & \new_Sorter100|11268_ ;
  assign \new_Sorter100|11368_  = \new_Sorter100|11267_  | \new_Sorter100|11268_ ;
  assign \new_Sorter100|11369_  = \new_Sorter100|11269_  & \new_Sorter100|11270_ ;
  assign \new_Sorter100|11370_  = \new_Sorter100|11269_  | \new_Sorter100|11270_ ;
  assign \new_Sorter100|11371_  = \new_Sorter100|11271_  & \new_Sorter100|11272_ ;
  assign \new_Sorter100|11372_  = \new_Sorter100|11271_  | \new_Sorter100|11272_ ;
  assign \new_Sorter100|11373_  = \new_Sorter100|11273_  & \new_Sorter100|11274_ ;
  assign \new_Sorter100|11374_  = \new_Sorter100|11273_  | \new_Sorter100|11274_ ;
  assign \new_Sorter100|11375_  = \new_Sorter100|11275_  & \new_Sorter100|11276_ ;
  assign \new_Sorter100|11376_  = \new_Sorter100|11275_  | \new_Sorter100|11276_ ;
  assign \new_Sorter100|11377_  = \new_Sorter100|11277_  & \new_Sorter100|11278_ ;
  assign \new_Sorter100|11378_  = \new_Sorter100|11277_  | \new_Sorter100|11278_ ;
  assign \new_Sorter100|11379_  = \new_Sorter100|11279_  & \new_Sorter100|11280_ ;
  assign \new_Sorter100|11380_  = \new_Sorter100|11279_  | \new_Sorter100|11280_ ;
  assign \new_Sorter100|11381_  = \new_Sorter100|11281_  & \new_Sorter100|11282_ ;
  assign \new_Sorter100|11382_  = \new_Sorter100|11281_  | \new_Sorter100|11282_ ;
  assign \new_Sorter100|11383_  = \new_Sorter100|11283_  & \new_Sorter100|11284_ ;
  assign \new_Sorter100|11384_  = \new_Sorter100|11283_  | \new_Sorter100|11284_ ;
  assign \new_Sorter100|11385_  = \new_Sorter100|11285_  & \new_Sorter100|11286_ ;
  assign \new_Sorter100|11386_  = \new_Sorter100|11285_  | \new_Sorter100|11286_ ;
  assign \new_Sorter100|11387_  = \new_Sorter100|11287_  & \new_Sorter100|11288_ ;
  assign \new_Sorter100|11388_  = \new_Sorter100|11287_  | \new_Sorter100|11288_ ;
  assign \new_Sorter100|11389_  = \new_Sorter100|11289_  & \new_Sorter100|11290_ ;
  assign \new_Sorter100|11390_  = \new_Sorter100|11289_  | \new_Sorter100|11290_ ;
  assign \new_Sorter100|11391_  = \new_Sorter100|11291_  & \new_Sorter100|11292_ ;
  assign \new_Sorter100|11392_  = \new_Sorter100|11291_  | \new_Sorter100|11292_ ;
  assign \new_Sorter100|11393_  = \new_Sorter100|11293_  & \new_Sorter100|11294_ ;
  assign \new_Sorter100|11394_  = \new_Sorter100|11293_  | \new_Sorter100|11294_ ;
  assign \new_Sorter100|11395_  = \new_Sorter100|11295_  & \new_Sorter100|11296_ ;
  assign \new_Sorter100|11396_  = \new_Sorter100|11295_  | \new_Sorter100|11296_ ;
  assign \new_Sorter100|11397_  = \new_Sorter100|11297_  & \new_Sorter100|11298_ ;
  assign \new_Sorter100|11398_  = \new_Sorter100|11297_  | \new_Sorter100|11298_ ;
  assign \new_Sorter100|11400_  = \new_Sorter100|11300_  & \new_Sorter100|11301_ ;
  assign \new_Sorter100|11401_  = \new_Sorter100|11300_  | \new_Sorter100|11301_ ;
  assign \new_Sorter100|11402_  = \new_Sorter100|11302_  & \new_Sorter100|11303_ ;
  assign \new_Sorter100|11403_  = \new_Sorter100|11302_  | \new_Sorter100|11303_ ;
  assign \new_Sorter100|11404_  = \new_Sorter100|11304_  & \new_Sorter100|11305_ ;
  assign \new_Sorter100|11405_  = \new_Sorter100|11304_  | \new_Sorter100|11305_ ;
  assign \new_Sorter100|11406_  = \new_Sorter100|11306_  & \new_Sorter100|11307_ ;
  assign \new_Sorter100|11407_  = \new_Sorter100|11306_  | \new_Sorter100|11307_ ;
  assign \new_Sorter100|11408_  = \new_Sorter100|11308_  & \new_Sorter100|11309_ ;
  assign \new_Sorter100|11409_  = \new_Sorter100|11308_  | \new_Sorter100|11309_ ;
  assign \new_Sorter100|11410_  = \new_Sorter100|11310_  & \new_Sorter100|11311_ ;
  assign \new_Sorter100|11411_  = \new_Sorter100|11310_  | \new_Sorter100|11311_ ;
  assign \new_Sorter100|11412_  = \new_Sorter100|11312_  & \new_Sorter100|11313_ ;
  assign \new_Sorter100|11413_  = \new_Sorter100|11312_  | \new_Sorter100|11313_ ;
  assign \new_Sorter100|11414_  = \new_Sorter100|11314_  & \new_Sorter100|11315_ ;
  assign \new_Sorter100|11415_  = \new_Sorter100|11314_  | \new_Sorter100|11315_ ;
  assign \new_Sorter100|11416_  = \new_Sorter100|11316_  & \new_Sorter100|11317_ ;
  assign \new_Sorter100|11417_  = \new_Sorter100|11316_  | \new_Sorter100|11317_ ;
  assign \new_Sorter100|11418_  = \new_Sorter100|11318_  & \new_Sorter100|11319_ ;
  assign \new_Sorter100|11419_  = \new_Sorter100|11318_  | \new_Sorter100|11319_ ;
  assign \new_Sorter100|11420_  = \new_Sorter100|11320_  & \new_Sorter100|11321_ ;
  assign \new_Sorter100|11421_  = \new_Sorter100|11320_  | \new_Sorter100|11321_ ;
  assign \new_Sorter100|11422_  = \new_Sorter100|11322_  & \new_Sorter100|11323_ ;
  assign \new_Sorter100|11423_  = \new_Sorter100|11322_  | \new_Sorter100|11323_ ;
  assign \new_Sorter100|11424_  = \new_Sorter100|11324_  & \new_Sorter100|11325_ ;
  assign \new_Sorter100|11425_  = \new_Sorter100|11324_  | \new_Sorter100|11325_ ;
  assign \new_Sorter100|11426_  = \new_Sorter100|11326_  & \new_Sorter100|11327_ ;
  assign \new_Sorter100|11427_  = \new_Sorter100|11326_  | \new_Sorter100|11327_ ;
  assign \new_Sorter100|11428_  = \new_Sorter100|11328_  & \new_Sorter100|11329_ ;
  assign \new_Sorter100|11429_  = \new_Sorter100|11328_  | \new_Sorter100|11329_ ;
  assign \new_Sorter100|11430_  = \new_Sorter100|11330_  & \new_Sorter100|11331_ ;
  assign \new_Sorter100|11431_  = \new_Sorter100|11330_  | \new_Sorter100|11331_ ;
  assign \new_Sorter100|11432_  = \new_Sorter100|11332_  & \new_Sorter100|11333_ ;
  assign \new_Sorter100|11433_  = \new_Sorter100|11332_  | \new_Sorter100|11333_ ;
  assign \new_Sorter100|11434_  = \new_Sorter100|11334_  & \new_Sorter100|11335_ ;
  assign \new_Sorter100|11435_  = \new_Sorter100|11334_  | \new_Sorter100|11335_ ;
  assign \new_Sorter100|11436_  = \new_Sorter100|11336_  & \new_Sorter100|11337_ ;
  assign \new_Sorter100|11437_  = \new_Sorter100|11336_  | \new_Sorter100|11337_ ;
  assign \new_Sorter100|11438_  = \new_Sorter100|11338_  & \new_Sorter100|11339_ ;
  assign \new_Sorter100|11439_  = \new_Sorter100|11338_  | \new_Sorter100|11339_ ;
  assign \new_Sorter100|11440_  = \new_Sorter100|11340_  & \new_Sorter100|11341_ ;
  assign \new_Sorter100|11441_  = \new_Sorter100|11340_  | \new_Sorter100|11341_ ;
  assign \new_Sorter100|11442_  = \new_Sorter100|11342_  & \new_Sorter100|11343_ ;
  assign \new_Sorter100|11443_  = \new_Sorter100|11342_  | \new_Sorter100|11343_ ;
  assign \new_Sorter100|11444_  = \new_Sorter100|11344_  & \new_Sorter100|11345_ ;
  assign \new_Sorter100|11445_  = \new_Sorter100|11344_  | \new_Sorter100|11345_ ;
  assign \new_Sorter100|11446_  = \new_Sorter100|11346_  & \new_Sorter100|11347_ ;
  assign \new_Sorter100|11447_  = \new_Sorter100|11346_  | \new_Sorter100|11347_ ;
  assign \new_Sorter100|11448_  = \new_Sorter100|11348_  & \new_Sorter100|11349_ ;
  assign \new_Sorter100|11449_  = \new_Sorter100|11348_  | \new_Sorter100|11349_ ;
  assign \new_Sorter100|11450_  = \new_Sorter100|11350_  & \new_Sorter100|11351_ ;
  assign \new_Sorter100|11451_  = \new_Sorter100|11350_  | \new_Sorter100|11351_ ;
  assign \new_Sorter100|11452_  = \new_Sorter100|11352_  & \new_Sorter100|11353_ ;
  assign \new_Sorter100|11453_  = \new_Sorter100|11352_  | \new_Sorter100|11353_ ;
  assign \new_Sorter100|11454_  = \new_Sorter100|11354_  & \new_Sorter100|11355_ ;
  assign \new_Sorter100|11455_  = \new_Sorter100|11354_  | \new_Sorter100|11355_ ;
  assign \new_Sorter100|11456_  = \new_Sorter100|11356_  & \new_Sorter100|11357_ ;
  assign \new_Sorter100|11457_  = \new_Sorter100|11356_  | \new_Sorter100|11357_ ;
  assign \new_Sorter100|11458_  = \new_Sorter100|11358_  & \new_Sorter100|11359_ ;
  assign \new_Sorter100|11459_  = \new_Sorter100|11358_  | \new_Sorter100|11359_ ;
  assign \new_Sorter100|11460_  = \new_Sorter100|11360_  & \new_Sorter100|11361_ ;
  assign \new_Sorter100|11461_  = \new_Sorter100|11360_  | \new_Sorter100|11361_ ;
  assign \new_Sorter100|11462_  = \new_Sorter100|11362_  & \new_Sorter100|11363_ ;
  assign \new_Sorter100|11463_  = \new_Sorter100|11362_  | \new_Sorter100|11363_ ;
  assign \new_Sorter100|11464_  = \new_Sorter100|11364_  & \new_Sorter100|11365_ ;
  assign \new_Sorter100|11465_  = \new_Sorter100|11364_  | \new_Sorter100|11365_ ;
  assign \new_Sorter100|11466_  = \new_Sorter100|11366_  & \new_Sorter100|11367_ ;
  assign \new_Sorter100|11467_  = \new_Sorter100|11366_  | \new_Sorter100|11367_ ;
  assign \new_Sorter100|11468_  = \new_Sorter100|11368_  & \new_Sorter100|11369_ ;
  assign \new_Sorter100|11469_  = \new_Sorter100|11368_  | \new_Sorter100|11369_ ;
  assign \new_Sorter100|11470_  = \new_Sorter100|11370_  & \new_Sorter100|11371_ ;
  assign \new_Sorter100|11471_  = \new_Sorter100|11370_  | \new_Sorter100|11371_ ;
  assign \new_Sorter100|11472_  = \new_Sorter100|11372_  & \new_Sorter100|11373_ ;
  assign \new_Sorter100|11473_  = \new_Sorter100|11372_  | \new_Sorter100|11373_ ;
  assign \new_Sorter100|11474_  = \new_Sorter100|11374_  & \new_Sorter100|11375_ ;
  assign \new_Sorter100|11475_  = \new_Sorter100|11374_  | \new_Sorter100|11375_ ;
  assign \new_Sorter100|11476_  = \new_Sorter100|11376_  & \new_Sorter100|11377_ ;
  assign \new_Sorter100|11477_  = \new_Sorter100|11376_  | \new_Sorter100|11377_ ;
  assign \new_Sorter100|11478_  = \new_Sorter100|11378_  & \new_Sorter100|11379_ ;
  assign \new_Sorter100|11479_  = \new_Sorter100|11378_  | \new_Sorter100|11379_ ;
  assign \new_Sorter100|11480_  = \new_Sorter100|11380_  & \new_Sorter100|11381_ ;
  assign \new_Sorter100|11481_  = \new_Sorter100|11380_  | \new_Sorter100|11381_ ;
  assign \new_Sorter100|11482_  = \new_Sorter100|11382_  & \new_Sorter100|11383_ ;
  assign \new_Sorter100|11483_  = \new_Sorter100|11382_  | \new_Sorter100|11383_ ;
  assign \new_Sorter100|11484_  = \new_Sorter100|11384_  & \new_Sorter100|11385_ ;
  assign \new_Sorter100|11485_  = \new_Sorter100|11384_  | \new_Sorter100|11385_ ;
  assign \new_Sorter100|11486_  = \new_Sorter100|11386_  & \new_Sorter100|11387_ ;
  assign \new_Sorter100|11487_  = \new_Sorter100|11386_  | \new_Sorter100|11387_ ;
  assign \new_Sorter100|11488_  = \new_Sorter100|11388_  & \new_Sorter100|11389_ ;
  assign \new_Sorter100|11489_  = \new_Sorter100|11388_  | \new_Sorter100|11389_ ;
  assign \new_Sorter100|11490_  = \new_Sorter100|11390_  & \new_Sorter100|11391_ ;
  assign \new_Sorter100|11491_  = \new_Sorter100|11390_  | \new_Sorter100|11391_ ;
  assign \new_Sorter100|11492_  = \new_Sorter100|11392_  & \new_Sorter100|11393_ ;
  assign \new_Sorter100|11493_  = \new_Sorter100|11392_  | \new_Sorter100|11393_ ;
  assign \new_Sorter100|11494_  = \new_Sorter100|11394_  & \new_Sorter100|11395_ ;
  assign \new_Sorter100|11495_  = \new_Sorter100|11394_  | \new_Sorter100|11395_ ;
  assign \new_Sorter100|11496_  = \new_Sorter100|11396_  & \new_Sorter100|11397_ ;
  assign \new_Sorter100|11497_  = \new_Sorter100|11396_  | \new_Sorter100|11397_ ;
  assign \new_Sorter100|11498_  = \new_Sorter100|11398_  & \new_Sorter100|11399_ ;
  assign \new_Sorter100|11499_  = \new_Sorter100|11398_  | \new_Sorter100|11399_ ;
  assign \new_Sorter100|11500_  = \new_Sorter100|11400_ ;
  assign \new_Sorter100|11599_  = \new_Sorter100|11499_ ;
  assign \new_Sorter100|11501_  = \new_Sorter100|11401_  & \new_Sorter100|11402_ ;
  assign \new_Sorter100|11502_  = \new_Sorter100|11401_  | \new_Sorter100|11402_ ;
  assign \new_Sorter100|11503_  = \new_Sorter100|11403_  & \new_Sorter100|11404_ ;
  assign \new_Sorter100|11504_  = \new_Sorter100|11403_  | \new_Sorter100|11404_ ;
  assign \new_Sorter100|11505_  = \new_Sorter100|11405_  & \new_Sorter100|11406_ ;
  assign \new_Sorter100|11506_  = \new_Sorter100|11405_  | \new_Sorter100|11406_ ;
  assign \new_Sorter100|11507_  = \new_Sorter100|11407_  & \new_Sorter100|11408_ ;
  assign \new_Sorter100|11508_  = \new_Sorter100|11407_  | \new_Sorter100|11408_ ;
  assign \new_Sorter100|11509_  = \new_Sorter100|11409_  & \new_Sorter100|11410_ ;
  assign \new_Sorter100|11510_  = \new_Sorter100|11409_  | \new_Sorter100|11410_ ;
  assign \new_Sorter100|11511_  = \new_Sorter100|11411_  & \new_Sorter100|11412_ ;
  assign \new_Sorter100|11512_  = \new_Sorter100|11411_  | \new_Sorter100|11412_ ;
  assign \new_Sorter100|11513_  = \new_Sorter100|11413_  & \new_Sorter100|11414_ ;
  assign \new_Sorter100|11514_  = \new_Sorter100|11413_  | \new_Sorter100|11414_ ;
  assign \new_Sorter100|11515_  = \new_Sorter100|11415_  & \new_Sorter100|11416_ ;
  assign \new_Sorter100|11516_  = \new_Sorter100|11415_  | \new_Sorter100|11416_ ;
  assign \new_Sorter100|11517_  = \new_Sorter100|11417_  & \new_Sorter100|11418_ ;
  assign \new_Sorter100|11518_  = \new_Sorter100|11417_  | \new_Sorter100|11418_ ;
  assign \new_Sorter100|11519_  = \new_Sorter100|11419_  & \new_Sorter100|11420_ ;
  assign \new_Sorter100|11520_  = \new_Sorter100|11419_  | \new_Sorter100|11420_ ;
  assign \new_Sorter100|11521_  = \new_Sorter100|11421_  & \new_Sorter100|11422_ ;
  assign \new_Sorter100|11522_  = \new_Sorter100|11421_  | \new_Sorter100|11422_ ;
  assign \new_Sorter100|11523_  = \new_Sorter100|11423_  & \new_Sorter100|11424_ ;
  assign \new_Sorter100|11524_  = \new_Sorter100|11423_  | \new_Sorter100|11424_ ;
  assign \new_Sorter100|11525_  = \new_Sorter100|11425_  & \new_Sorter100|11426_ ;
  assign \new_Sorter100|11526_  = \new_Sorter100|11425_  | \new_Sorter100|11426_ ;
  assign \new_Sorter100|11527_  = \new_Sorter100|11427_  & \new_Sorter100|11428_ ;
  assign \new_Sorter100|11528_  = \new_Sorter100|11427_  | \new_Sorter100|11428_ ;
  assign \new_Sorter100|11529_  = \new_Sorter100|11429_  & \new_Sorter100|11430_ ;
  assign \new_Sorter100|11530_  = \new_Sorter100|11429_  | \new_Sorter100|11430_ ;
  assign \new_Sorter100|11531_  = \new_Sorter100|11431_  & \new_Sorter100|11432_ ;
  assign \new_Sorter100|11532_  = \new_Sorter100|11431_  | \new_Sorter100|11432_ ;
  assign \new_Sorter100|11533_  = \new_Sorter100|11433_  & \new_Sorter100|11434_ ;
  assign \new_Sorter100|11534_  = \new_Sorter100|11433_  | \new_Sorter100|11434_ ;
  assign \new_Sorter100|11535_  = \new_Sorter100|11435_  & \new_Sorter100|11436_ ;
  assign \new_Sorter100|11536_  = \new_Sorter100|11435_  | \new_Sorter100|11436_ ;
  assign \new_Sorter100|11537_  = \new_Sorter100|11437_  & \new_Sorter100|11438_ ;
  assign \new_Sorter100|11538_  = \new_Sorter100|11437_  | \new_Sorter100|11438_ ;
  assign \new_Sorter100|11539_  = \new_Sorter100|11439_  & \new_Sorter100|11440_ ;
  assign \new_Sorter100|11540_  = \new_Sorter100|11439_  | \new_Sorter100|11440_ ;
  assign \new_Sorter100|11541_  = \new_Sorter100|11441_  & \new_Sorter100|11442_ ;
  assign \new_Sorter100|11542_  = \new_Sorter100|11441_  | \new_Sorter100|11442_ ;
  assign \new_Sorter100|11543_  = \new_Sorter100|11443_  & \new_Sorter100|11444_ ;
  assign \new_Sorter100|11544_  = \new_Sorter100|11443_  | \new_Sorter100|11444_ ;
  assign \new_Sorter100|11545_  = \new_Sorter100|11445_  & \new_Sorter100|11446_ ;
  assign \new_Sorter100|11546_  = \new_Sorter100|11445_  | \new_Sorter100|11446_ ;
  assign \new_Sorter100|11547_  = \new_Sorter100|11447_  & \new_Sorter100|11448_ ;
  assign \new_Sorter100|11548_  = \new_Sorter100|11447_  | \new_Sorter100|11448_ ;
  assign \new_Sorter100|11549_  = \new_Sorter100|11449_  & \new_Sorter100|11450_ ;
  assign \new_Sorter100|11550_  = \new_Sorter100|11449_  | \new_Sorter100|11450_ ;
  assign \new_Sorter100|11551_  = \new_Sorter100|11451_  & \new_Sorter100|11452_ ;
  assign \new_Sorter100|11552_  = \new_Sorter100|11451_  | \new_Sorter100|11452_ ;
  assign \new_Sorter100|11553_  = \new_Sorter100|11453_  & \new_Sorter100|11454_ ;
  assign \new_Sorter100|11554_  = \new_Sorter100|11453_  | \new_Sorter100|11454_ ;
  assign \new_Sorter100|11555_  = \new_Sorter100|11455_  & \new_Sorter100|11456_ ;
  assign \new_Sorter100|11556_  = \new_Sorter100|11455_  | \new_Sorter100|11456_ ;
  assign \new_Sorter100|11557_  = \new_Sorter100|11457_  & \new_Sorter100|11458_ ;
  assign \new_Sorter100|11558_  = \new_Sorter100|11457_  | \new_Sorter100|11458_ ;
  assign \new_Sorter100|11559_  = \new_Sorter100|11459_  & \new_Sorter100|11460_ ;
  assign \new_Sorter100|11560_  = \new_Sorter100|11459_  | \new_Sorter100|11460_ ;
  assign \new_Sorter100|11561_  = \new_Sorter100|11461_  & \new_Sorter100|11462_ ;
  assign \new_Sorter100|11562_  = \new_Sorter100|11461_  | \new_Sorter100|11462_ ;
  assign \new_Sorter100|11563_  = \new_Sorter100|11463_  & \new_Sorter100|11464_ ;
  assign \new_Sorter100|11564_  = \new_Sorter100|11463_  | \new_Sorter100|11464_ ;
  assign \new_Sorter100|11565_  = \new_Sorter100|11465_  & \new_Sorter100|11466_ ;
  assign \new_Sorter100|11566_  = \new_Sorter100|11465_  | \new_Sorter100|11466_ ;
  assign \new_Sorter100|11567_  = \new_Sorter100|11467_  & \new_Sorter100|11468_ ;
  assign \new_Sorter100|11568_  = \new_Sorter100|11467_  | \new_Sorter100|11468_ ;
  assign \new_Sorter100|11569_  = \new_Sorter100|11469_  & \new_Sorter100|11470_ ;
  assign \new_Sorter100|11570_  = \new_Sorter100|11469_  | \new_Sorter100|11470_ ;
  assign \new_Sorter100|11571_  = \new_Sorter100|11471_  & \new_Sorter100|11472_ ;
  assign \new_Sorter100|11572_  = \new_Sorter100|11471_  | \new_Sorter100|11472_ ;
  assign \new_Sorter100|11573_  = \new_Sorter100|11473_  & \new_Sorter100|11474_ ;
  assign \new_Sorter100|11574_  = \new_Sorter100|11473_  | \new_Sorter100|11474_ ;
  assign \new_Sorter100|11575_  = \new_Sorter100|11475_  & \new_Sorter100|11476_ ;
  assign \new_Sorter100|11576_  = \new_Sorter100|11475_  | \new_Sorter100|11476_ ;
  assign \new_Sorter100|11577_  = \new_Sorter100|11477_  & \new_Sorter100|11478_ ;
  assign \new_Sorter100|11578_  = \new_Sorter100|11477_  | \new_Sorter100|11478_ ;
  assign \new_Sorter100|11579_  = \new_Sorter100|11479_  & \new_Sorter100|11480_ ;
  assign \new_Sorter100|11580_  = \new_Sorter100|11479_  | \new_Sorter100|11480_ ;
  assign \new_Sorter100|11581_  = \new_Sorter100|11481_  & \new_Sorter100|11482_ ;
  assign \new_Sorter100|11582_  = \new_Sorter100|11481_  | \new_Sorter100|11482_ ;
  assign \new_Sorter100|11583_  = \new_Sorter100|11483_  & \new_Sorter100|11484_ ;
  assign \new_Sorter100|11584_  = \new_Sorter100|11483_  | \new_Sorter100|11484_ ;
  assign \new_Sorter100|11585_  = \new_Sorter100|11485_  & \new_Sorter100|11486_ ;
  assign \new_Sorter100|11586_  = \new_Sorter100|11485_  | \new_Sorter100|11486_ ;
  assign \new_Sorter100|11587_  = \new_Sorter100|11487_  & \new_Sorter100|11488_ ;
  assign \new_Sorter100|11588_  = \new_Sorter100|11487_  | \new_Sorter100|11488_ ;
  assign \new_Sorter100|11589_  = \new_Sorter100|11489_  & \new_Sorter100|11490_ ;
  assign \new_Sorter100|11590_  = \new_Sorter100|11489_  | \new_Sorter100|11490_ ;
  assign \new_Sorter100|11591_  = \new_Sorter100|11491_  & \new_Sorter100|11492_ ;
  assign \new_Sorter100|11592_  = \new_Sorter100|11491_  | \new_Sorter100|11492_ ;
  assign \new_Sorter100|11593_  = \new_Sorter100|11493_  & \new_Sorter100|11494_ ;
  assign \new_Sorter100|11594_  = \new_Sorter100|11493_  | \new_Sorter100|11494_ ;
  assign \new_Sorter100|11595_  = \new_Sorter100|11495_  & \new_Sorter100|11496_ ;
  assign \new_Sorter100|11596_  = \new_Sorter100|11495_  | \new_Sorter100|11496_ ;
  assign \new_Sorter100|11597_  = \new_Sorter100|11497_  & \new_Sorter100|11498_ ;
  assign \new_Sorter100|11598_  = \new_Sorter100|11497_  | \new_Sorter100|11498_ ;
  assign \new_Sorter100|11600_  = \new_Sorter100|11500_  & \new_Sorter100|11501_ ;
  assign \new_Sorter100|11601_  = \new_Sorter100|11500_  | \new_Sorter100|11501_ ;
  assign \new_Sorter100|11602_  = \new_Sorter100|11502_  & \new_Sorter100|11503_ ;
  assign \new_Sorter100|11603_  = \new_Sorter100|11502_  | \new_Sorter100|11503_ ;
  assign \new_Sorter100|11604_  = \new_Sorter100|11504_  & \new_Sorter100|11505_ ;
  assign \new_Sorter100|11605_  = \new_Sorter100|11504_  | \new_Sorter100|11505_ ;
  assign \new_Sorter100|11606_  = \new_Sorter100|11506_  & \new_Sorter100|11507_ ;
  assign \new_Sorter100|11607_  = \new_Sorter100|11506_  | \new_Sorter100|11507_ ;
  assign \new_Sorter100|11608_  = \new_Sorter100|11508_  & \new_Sorter100|11509_ ;
  assign \new_Sorter100|11609_  = \new_Sorter100|11508_  | \new_Sorter100|11509_ ;
  assign \new_Sorter100|11610_  = \new_Sorter100|11510_  & \new_Sorter100|11511_ ;
  assign \new_Sorter100|11611_  = \new_Sorter100|11510_  | \new_Sorter100|11511_ ;
  assign \new_Sorter100|11612_  = \new_Sorter100|11512_  & \new_Sorter100|11513_ ;
  assign \new_Sorter100|11613_  = \new_Sorter100|11512_  | \new_Sorter100|11513_ ;
  assign \new_Sorter100|11614_  = \new_Sorter100|11514_  & \new_Sorter100|11515_ ;
  assign \new_Sorter100|11615_  = \new_Sorter100|11514_  | \new_Sorter100|11515_ ;
  assign \new_Sorter100|11616_  = \new_Sorter100|11516_  & \new_Sorter100|11517_ ;
  assign \new_Sorter100|11617_  = \new_Sorter100|11516_  | \new_Sorter100|11517_ ;
  assign \new_Sorter100|11618_  = \new_Sorter100|11518_  & \new_Sorter100|11519_ ;
  assign \new_Sorter100|11619_  = \new_Sorter100|11518_  | \new_Sorter100|11519_ ;
  assign \new_Sorter100|11620_  = \new_Sorter100|11520_  & \new_Sorter100|11521_ ;
  assign \new_Sorter100|11621_  = \new_Sorter100|11520_  | \new_Sorter100|11521_ ;
  assign \new_Sorter100|11622_  = \new_Sorter100|11522_  & \new_Sorter100|11523_ ;
  assign \new_Sorter100|11623_  = \new_Sorter100|11522_  | \new_Sorter100|11523_ ;
  assign \new_Sorter100|11624_  = \new_Sorter100|11524_  & \new_Sorter100|11525_ ;
  assign \new_Sorter100|11625_  = \new_Sorter100|11524_  | \new_Sorter100|11525_ ;
  assign \new_Sorter100|11626_  = \new_Sorter100|11526_  & \new_Sorter100|11527_ ;
  assign \new_Sorter100|11627_  = \new_Sorter100|11526_  | \new_Sorter100|11527_ ;
  assign \new_Sorter100|11628_  = \new_Sorter100|11528_  & \new_Sorter100|11529_ ;
  assign \new_Sorter100|11629_  = \new_Sorter100|11528_  | \new_Sorter100|11529_ ;
  assign \new_Sorter100|11630_  = \new_Sorter100|11530_  & \new_Sorter100|11531_ ;
  assign \new_Sorter100|11631_  = \new_Sorter100|11530_  | \new_Sorter100|11531_ ;
  assign \new_Sorter100|11632_  = \new_Sorter100|11532_  & \new_Sorter100|11533_ ;
  assign \new_Sorter100|11633_  = \new_Sorter100|11532_  | \new_Sorter100|11533_ ;
  assign \new_Sorter100|11634_  = \new_Sorter100|11534_  & \new_Sorter100|11535_ ;
  assign \new_Sorter100|11635_  = \new_Sorter100|11534_  | \new_Sorter100|11535_ ;
  assign \new_Sorter100|11636_  = \new_Sorter100|11536_  & \new_Sorter100|11537_ ;
  assign \new_Sorter100|11637_  = \new_Sorter100|11536_  | \new_Sorter100|11537_ ;
  assign \new_Sorter100|11638_  = \new_Sorter100|11538_  & \new_Sorter100|11539_ ;
  assign \new_Sorter100|11639_  = \new_Sorter100|11538_  | \new_Sorter100|11539_ ;
  assign \new_Sorter100|11640_  = \new_Sorter100|11540_  & \new_Sorter100|11541_ ;
  assign \new_Sorter100|11641_  = \new_Sorter100|11540_  | \new_Sorter100|11541_ ;
  assign \new_Sorter100|11642_  = \new_Sorter100|11542_  & \new_Sorter100|11543_ ;
  assign \new_Sorter100|11643_  = \new_Sorter100|11542_  | \new_Sorter100|11543_ ;
  assign \new_Sorter100|11644_  = \new_Sorter100|11544_  & \new_Sorter100|11545_ ;
  assign \new_Sorter100|11645_  = \new_Sorter100|11544_  | \new_Sorter100|11545_ ;
  assign \new_Sorter100|11646_  = \new_Sorter100|11546_  & \new_Sorter100|11547_ ;
  assign \new_Sorter100|11647_  = \new_Sorter100|11546_  | \new_Sorter100|11547_ ;
  assign \new_Sorter100|11648_  = \new_Sorter100|11548_  & \new_Sorter100|11549_ ;
  assign \new_Sorter100|11649_  = \new_Sorter100|11548_  | \new_Sorter100|11549_ ;
  assign \new_Sorter100|11650_  = \new_Sorter100|11550_  & \new_Sorter100|11551_ ;
  assign \new_Sorter100|11651_  = \new_Sorter100|11550_  | \new_Sorter100|11551_ ;
  assign \new_Sorter100|11652_  = \new_Sorter100|11552_  & \new_Sorter100|11553_ ;
  assign \new_Sorter100|11653_  = \new_Sorter100|11552_  | \new_Sorter100|11553_ ;
  assign \new_Sorter100|11654_  = \new_Sorter100|11554_  & \new_Sorter100|11555_ ;
  assign \new_Sorter100|11655_  = \new_Sorter100|11554_  | \new_Sorter100|11555_ ;
  assign \new_Sorter100|11656_  = \new_Sorter100|11556_  & \new_Sorter100|11557_ ;
  assign \new_Sorter100|11657_  = \new_Sorter100|11556_  | \new_Sorter100|11557_ ;
  assign \new_Sorter100|11658_  = \new_Sorter100|11558_  & \new_Sorter100|11559_ ;
  assign \new_Sorter100|11659_  = \new_Sorter100|11558_  | \new_Sorter100|11559_ ;
  assign \new_Sorter100|11660_  = \new_Sorter100|11560_  & \new_Sorter100|11561_ ;
  assign \new_Sorter100|11661_  = \new_Sorter100|11560_  | \new_Sorter100|11561_ ;
  assign \new_Sorter100|11662_  = \new_Sorter100|11562_  & \new_Sorter100|11563_ ;
  assign \new_Sorter100|11663_  = \new_Sorter100|11562_  | \new_Sorter100|11563_ ;
  assign \new_Sorter100|11664_  = \new_Sorter100|11564_  & \new_Sorter100|11565_ ;
  assign \new_Sorter100|11665_  = \new_Sorter100|11564_  | \new_Sorter100|11565_ ;
  assign \new_Sorter100|11666_  = \new_Sorter100|11566_  & \new_Sorter100|11567_ ;
  assign \new_Sorter100|11667_  = \new_Sorter100|11566_  | \new_Sorter100|11567_ ;
  assign \new_Sorter100|11668_  = \new_Sorter100|11568_  & \new_Sorter100|11569_ ;
  assign \new_Sorter100|11669_  = \new_Sorter100|11568_  | \new_Sorter100|11569_ ;
  assign \new_Sorter100|11670_  = \new_Sorter100|11570_  & \new_Sorter100|11571_ ;
  assign \new_Sorter100|11671_  = \new_Sorter100|11570_  | \new_Sorter100|11571_ ;
  assign \new_Sorter100|11672_  = \new_Sorter100|11572_  & \new_Sorter100|11573_ ;
  assign \new_Sorter100|11673_  = \new_Sorter100|11572_  | \new_Sorter100|11573_ ;
  assign \new_Sorter100|11674_  = \new_Sorter100|11574_  & \new_Sorter100|11575_ ;
  assign \new_Sorter100|11675_  = \new_Sorter100|11574_  | \new_Sorter100|11575_ ;
  assign \new_Sorter100|11676_  = \new_Sorter100|11576_  & \new_Sorter100|11577_ ;
  assign \new_Sorter100|11677_  = \new_Sorter100|11576_  | \new_Sorter100|11577_ ;
  assign \new_Sorter100|11678_  = \new_Sorter100|11578_  & \new_Sorter100|11579_ ;
  assign \new_Sorter100|11679_  = \new_Sorter100|11578_  | \new_Sorter100|11579_ ;
  assign \new_Sorter100|11680_  = \new_Sorter100|11580_  & \new_Sorter100|11581_ ;
  assign \new_Sorter100|11681_  = \new_Sorter100|11580_  | \new_Sorter100|11581_ ;
  assign \new_Sorter100|11682_  = \new_Sorter100|11582_  & \new_Sorter100|11583_ ;
  assign \new_Sorter100|11683_  = \new_Sorter100|11582_  | \new_Sorter100|11583_ ;
  assign \new_Sorter100|11684_  = \new_Sorter100|11584_  & \new_Sorter100|11585_ ;
  assign \new_Sorter100|11685_  = \new_Sorter100|11584_  | \new_Sorter100|11585_ ;
  assign \new_Sorter100|11686_  = \new_Sorter100|11586_  & \new_Sorter100|11587_ ;
  assign \new_Sorter100|11687_  = \new_Sorter100|11586_  | \new_Sorter100|11587_ ;
  assign \new_Sorter100|11688_  = \new_Sorter100|11588_  & \new_Sorter100|11589_ ;
  assign \new_Sorter100|11689_  = \new_Sorter100|11588_  | \new_Sorter100|11589_ ;
  assign \new_Sorter100|11690_  = \new_Sorter100|11590_  & \new_Sorter100|11591_ ;
  assign \new_Sorter100|11691_  = \new_Sorter100|11590_  | \new_Sorter100|11591_ ;
  assign \new_Sorter100|11692_  = \new_Sorter100|11592_  & \new_Sorter100|11593_ ;
  assign \new_Sorter100|11693_  = \new_Sorter100|11592_  | \new_Sorter100|11593_ ;
  assign \new_Sorter100|11694_  = \new_Sorter100|11594_  & \new_Sorter100|11595_ ;
  assign \new_Sorter100|11695_  = \new_Sorter100|11594_  | \new_Sorter100|11595_ ;
  assign \new_Sorter100|11696_  = \new_Sorter100|11596_  & \new_Sorter100|11597_ ;
  assign \new_Sorter100|11697_  = \new_Sorter100|11596_  | \new_Sorter100|11597_ ;
  assign \new_Sorter100|11698_  = \new_Sorter100|11598_  & \new_Sorter100|11599_ ;
  assign \new_Sorter100|11699_  = \new_Sorter100|11598_  | \new_Sorter100|11599_ ;
  assign \new_Sorter100|11700_  = \new_Sorter100|11600_ ;
  assign \new_Sorter100|11799_  = \new_Sorter100|11699_ ;
  assign \new_Sorter100|11701_  = \new_Sorter100|11601_  & \new_Sorter100|11602_ ;
  assign \new_Sorter100|11702_  = \new_Sorter100|11601_  | \new_Sorter100|11602_ ;
  assign \new_Sorter100|11703_  = \new_Sorter100|11603_  & \new_Sorter100|11604_ ;
  assign \new_Sorter100|11704_  = \new_Sorter100|11603_  | \new_Sorter100|11604_ ;
  assign \new_Sorter100|11705_  = \new_Sorter100|11605_  & \new_Sorter100|11606_ ;
  assign \new_Sorter100|11706_  = \new_Sorter100|11605_  | \new_Sorter100|11606_ ;
  assign \new_Sorter100|11707_  = \new_Sorter100|11607_  & \new_Sorter100|11608_ ;
  assign \new_Sorter100|11708_  = \new_Sorter100|11607_  | \new_Sorter100|11608_ ;
  assign \new_Sorter100|11709_  = \new_Sorter100|11609_  & \new_Sorter100|11610_ ;
  assign \new_Sorter100|11710_  = \new_Sorter100|11609_  | \new_Sorter100|11610_ ;
  assign \new_Sorter100|11711_  = \new_Sorter100|11611_  & \new_Sorter100|11612_ ;
  assign \new_Sorter100|11712_  = \new_Sorter100|11611_  | \new_Sorter100|11612_ ;
  assign \new_Sorter100|11713_  = \new_Sorter100|11613_  & \new_Sorter100|11614_ ;
  assign \new_Sorter100|11714_  = \new_Sorter100|11613_  | \new_Sorter100|11614_ ;
  assign \new_Sorter100|11715_  = \new_Sorter100|11615_  & \new_Sorter100|11616_ ;
  assign \new_Sorter100|11716_  = \new_Sorter100|11615_  | \new_Sorter100|11616_ ;
  assign \new_Sorter100|11717_  = \new_Sorter100|11617_  & \new_Sorter100|11618_ ;
  assign \new_Sorter100|11718_  = \new_Sorter100|11617_  | \new_Sorter100|11618_ ;
  assign \new_Sorter100|11719_  = \new_Sorter100|11619_  & \new_Sorter100|11620_ ;
  assign \new_Sorter100|11720_  = \new_Sorter100|11619_  | \new_Sorter100|11620_ ;
  assign \new_Sorter100|11721_  = \new_Sorter100|11621_  & \new_Sorter100|11622_ ;
  assign \new_Sorter100|11722_  = \new_Sorter100|11621_  | \new_Sorter100|11622_ ;
  assign \new_Sorter100|11723_  = \new_Sorter100|11623_  & \new_Sorter100|11624_ ;
  assign \new_Sorter100|11724_  = \new_Sorter100|11623_  | \new_Sorter100|11624_ ;
  assign \new_Sorter100|11725_  = \new_Sorter100|11625_  & \new_Sorter100|11626_ ;
  assign \new_Sorter100|11726_  = \new_Sorter100|11625_  | \new_Sorter100|11626_ ;
  assign \new_Sorter100|11727_  = \new_Sorter100|11627_  & \new_Sorter100|11628_ ;
  assign \new_Sorter100|11728_  = \new_Sorter100|11627_  | \new_Sorter100|11628_ ;
  assign \new_Sorter100|11729_  = \new_Sorter100|11629_  & \new_Sorter100|11630_ ;
  assign \new_Sorter100|11730_  = \new_Sorter100|11629_  | \new_Sorter100|11630_ ;
  assign \new_Sorter100|11731_  = \new_Sorter100|11631_  & \new_Sorter100|11632_ ;
  assign \new_Sorter100|11732_  = \new_Sorter100|11631_  | \new_Sorter100|11632_ ;
  assign \new_Sorter100|11733_  = \new_Sorter100|11633_  & \new_Sorter100|11634_ ;
  assign \new_Sorter100|11734_  = \new_Sorter100|11633_  | \new_Sorter100|11634_ ;
  assign \new_Sorter100|11735_  = \new_Sorter100|11635_  & \new_Sorter100|11636_ ;
  assign \new_Sorter100|11736_  = \new_Sorter100|11635_  | \new_Sorter100|11636_ ;
  assign \new_Sorter100|11737_  = \new_Sorter100|11637_  & \new_Sorter100|11638_ ;
  assign \new_Sorter100|11738_  = \new_Sorter100|11637_  | \new_Sorter100|11638_ ;
  assign \new_Sorter100|11739_  = \new_Sorter100|11639_  & \new_Sorter100|11640_ ;
  assign \new_Sorter100|11740_  = \new_Sorter100|11639_  | \new_Sorter100|11640_ ;
  assign \new_Sorter100|11741_  = \new_Sorter100|11641_  & \new_Sorter100|11642_ ;
  assign \new_Sorter100|11742_  = \new_Sorter100|11641_  | \new_Sorter100|11642_ ;
  assign \new_Sorter100|11743_  = \new_Sorter100|11643_  & \new_Sorter100|11644_ ;
  assign \new_Sorter100|11744_  = \new_Sorter100|11643_  | \new_Sorter100|11644_ ;
  assign \new_Sorter100|11745_  = \new_Sorter100|11645_  & \new_Sorter100|11646_ ;
  assign \new_Sorter100|11746_  = \new_Sorter100|11645_  | \new_Sorter100|11646_ ;
  assign \new_Sorter100|11747_  = \new_Sorter100|11647_  & \new_Sorter100|11648_ ;
  assign \new_Sorter100|11748_  = \new_Sorter100|11647_  | \new_Sorter100|11648_ ;
  assign \new_Sorter100|11749_  = \new_Sorter100|11649_  & \new_Sorter100|11650_ ;
  assign \new_Sorter100|11750_  = \new_Sorter100|11649_  | \new_Sorter100|11650_ ;
  assign \new_Sorter100|11751_  = \new_Sorter100|11651_  & \new_Sorter100|11652_ ;
  assign \new_Sorter100|11752_  = \new_Sorter100|11651_  | \new_Sorter100|11652_ ;
  assign \new_Sorter100|11753_  = \new_Sorter100|11653_  & \new_Sorter100|11654_ ;
  assign \new_Sorter100|11754_  = \new_Sorter100|11653_  | \new_Sorter100|11654_ ;
  assign \new_Sorter100|11755_  = \new_Sorter100|11655_  & \new_Sorter100|11656_ ;
  assign \new_Sorter100|11756_  = \new_Sorter100|11655_  | \new_Sorter100|11656_ ;
  assign \new_Sorter100|11757_  = \new_Sorter100|11657_  & \new_Sorter100|11658_ ;
  assign \new_Sorter100|11758_  = \new_Sorter100|11657_  | \new_Sorter100|11658_ ;
  assign \new_Sorter100|11759_  = \new_Sorter100|11659_  & \new_Sorter100|11660_ ;
  assign \new_Sorter100|11760_  = \new_Sorter100|11659_  | \new_Sorter100|11660_ ;
  assign \new_Sorter100|11761_  = \new_Sorter100|11661_  & \new_Sorter100|11662_ ;
  assign \new_Sorter100|11762_  = \new_Sorter100|11661_  | \new_Sorter100|11662_ ;
  assign \new_Sorter100|11763_  = \new_Sorter100|11663_  & \new_Sorter100|11664_ ;
  assign \new_Sorter100|11764_  = \new_Sorter100|11663_  | \new_Sorter100|11664_ ;
  assign \new_Sorter100|11765_  = \new_Sorter100|11665_  & \new_Sorter100|11666_ ;
  assign \new_Sorter100|11766_  = \new_Sorter100|11665_  | \new_Sorter100|11666_ ;
  assign \new_Sorter100|11767_  = \new_Sorter100|11667_  & \new_Sorter100|11668_ ;
  assign \new_Sorter100|11768_  = \new_Sorter100|11667_  | \new_Sorter100|11668_ ;
  assign \new_Sorter100|11769_  = \new_Sorter100|11669_  & \new_Sorter100|11670_ ;
  assign \new_Sorter100|11770_  = \new_Sorter100|11669_  | \new_Sorter100|11670_ ;
  assign \new_Sorter100|11771_  = \new_Sorter100|11671_  & \new_Sorter100|11672_ ;
  assign \new_Sorter100|11772_  = \new_Sorter100|11671_  | \new_Sorter100|11672_ ;
  assign \new_Sorter100|11773_  = \new_Sorter100|11673_  & \new_Sorter100|11674_ ;
  assign \new_Sorter100|11774_  = \new_Sorter100|11673_  | \new_Sorter100|11674_ ;
  assign \new_Sorter100|11775_  = \new_Sorter100|11675_  & \new_Sorter100|11676_ ;
  assign \new_Sorter100|11776_  = \new_Sorter100|11675_  | \new_Sorter100|11676_ ;
  assign \new_Sorter100|11777_  = \new_Sorter100|11677_  & \new_Sorter100|11678_ ;
  assign \new_Sorter100|11778_  = \new_Sorter100|11677_  | \new_Sorter100|11678_ ;
  assign \new_Sorter100|11779_  = \new_Sorter100|11679_  & \new_Sorter100|11680_ ;
  assign \new_Sorter100|11780_  = \new_Sorter100|11679_  | \new_Sorter100|11680_ ;
  assign \new_Sorter100|11781_  = \new_Sorter100|11681_  & \new_Sorter100|11682_ ;
  assign \new_Sorter100|11782_  = \new_Sorter100|11681_  | \new_Sorter100|11682_ ;
  assign \new_Sorter100|11783_  = \new_Sorter100|11683_  & \new_Sorter100|11684_ ;
  assign \new_Sorter100|11784_  = \new_Sorter100|11683_  | \new_Sorter100|11684_ ;
  assign \new_Sorter100|11785_  = \new_Sorter100|11685_  & \new_Sorter100|11686_ ;
  assign \new_Sorter100|11786_  = \new_Sorter100|11685_  | \new_Sorter100|11686_ ;
  assign \new_Sorter100|11787_  = \new_Sorter100|11687_  & \new_Sorter100|11688_ ;
  assign \new_Sorter100|11788_  = \new_Sorter100|11687_  | \new_Sorter100|11688_ ;
  assign \new_Sorter100|11789_  = \new_Sorter100|11689_  & \new_Sorter100|11690_ ;
  assign \new_Sorter100|11790_  = \new_Sorter100|11689_  | \new_Sorter100|11690_ ;
  assign \new_Sorter100|11791_  = \new_Sorter100|11691_  & \new_Sorter100|11692_ ;
  assign \new_Sorter100|11792_  = \new_Sorter100|11691_  | \new_Sorter100|11692_ ;
  assign \new_Sorter100|11793_  = \new_Sorter100|11693_  & \new_Sorter100|11694_ ;
  assign \new_Sorter100|11794_  = \new_Sorter100|11693_  | \new_Sorter100|11694_ ;
  assign \new_Sorter100|11795_  = \new_Sorter100|11695_  & \new_Sorter100|11696_ ;
  assign \new_Sorter100|11796_  = \new_Sorter100|11695_  | \new_Sorter100|11696_ ;
  assign \new_Sorter100|11797_  = \new_Sorter100|11697_  & \new_Sorter100|11698_ ;
  assign \new_Sorter100|11798_  = \new_Sorter100|11697_  | \new_Sorter100|11698_ ;
  assign \new_Sorter100|11800_  = \new_Sorter100|11700_  & \new_Sorter100|11701_ ;
  assign \new_Sorter100|11801_  = \new_Sorter100|11700_  | \new_Sorter100|11701_ ;
  assign \new_Sorter100|11802_  = \new_Sorter100|11702_  & \new_Sorter100|11703_ ;
  assign \new_Sorter100|11803_  = \new_Sorter100|11702_  | \new_Sorter100|11703_ ;
  assign \new_Sorter100|11804_  = \new_Sorter100|11704_  & \new_Sorter100|11705_ ;
  assign \new_Sorter100|11805_  = \new_Sorter100|11704_  | \new_Sorter100|11705_ ;
  assign \new_Sorter100|11806_  = \new_Sorter100|11706_  & \new_Sorter100|11707_ ;
  assign \new_Sorter100|11807_  = \new_Sorter100|11706_  | \new_Sorter100|11707_ ;
  assign \new_Sorter100|11808_  = \new_Sorter100|11708_  & \new_Sorter100|11709_ ;
  assign \new_Sorter100|11809_  = \new_Sorter100|11708_  | \new_Sorter100|11709_ ;
  assign \new_Sorter100|11810_  = \new_Sorter100|11710_  & \new_Sorter100|11711_ ;
  assign \new_Sorter100|11811_  = \new_Sorter100|11710_  | \new_Sorter100|11711_ ;
  assign \new_Sorter100|11812_  = \new_Sorter100|11712_  & \new_Sorter100|11713_ ;
  assign \new_Sorter100|11813_  = \new_Sorter100|11712_  | \new_Sorter100|11713_ ;
  assign \new_Sorter100|11814_  = \new_Sorter100|11714_  & \new_Sorter100|11715_ ;
  assign \new_Sorter100|11815_  = \new_Sorter100|11714_  | \new_Sorter100|11715_ ;
  assign \new_Sorter100|11816_  = \new_Sorter100|11716_  & \new_Sorter100|11717_ ;
  assign \new_Sorter100|11817_  = \new_Sorter100|11716_  | \new_Sorter100|11717_ ;
  assign \new_Sorter100|11818_  = \new_Sorter100|11718_  & \new_Sorter100|11719_ ;
  assign \new_Sorter100|11819_  = \new_Sorter100|11718_  | \new_Sorter100|11719_ ;
  assign \new_Sorter100|11820_  = \new_Sorter100|11720_  & \new_Sorter100|11721_ ;
  assign \new_Sorter100|11821_  = \new_Sorter100|11720_  | \new_Sorter100|11721_ ;
  assign \new_Sorter100|11822_  = \new_Sorter100|11722_  & \new_Sorter100|11723_ ;
  assign \new_Sorter100|11823_  = \new_Sorter100|11722_  | \new_Sorter100|11723_ ;
  assign \new_Sorter100|11824_  = \new_Sorter100|11724_  & \new_Sorter100|11725_ ;
  assign \new_Sorter100|11825_  = \new_Sorter100|11724_  | \new_Sorter100|11725_ ;
  assign \new_Sorter100|11826_  = \new_Sorter100|11726_  & \new_Sorter100|11727_ ;
  assign \new_Sorter100|11827_  = \new_Sorter100|11726_  | \new_Sorter100|11727_ ;
  assign \new_Sorter100|11828_  = \new_Sorter100|11728_  & \new_Sorter100|11729_ ;
  assign \new_Sorter100|11829_  = \new_Sorter100|11728_  | \new_Sorter100|11729_ ;
  assign \new_Sorter100|11830_  = \new_Sorter100|11730_  & \new_Sorter100|11731_ ;
  assign \new_Sorter100|11831_  = \new_Sorter100|11730_  | \new_Sorter100|11731_ ;
  assign \new_Sorter100|11832_  = \new_Sorter100|11732_  & \new_Sorter100|11733_ ;
  assign \new_Sorter100|11833_  = \new_Sorter100|11732_  | \new_Sorter100|11733_ ;
  assign \new_Sorter100|11834_  = \new_Sorter100|11734_  & \new_Sorter100|11735_ ;
  assign \new_Sorter100|11835_  = \new_Sorter100|11734_  | \new_Sorter100|11735_ ;
  assign \new_Sorter100|11836_  = \new_Sorter100|11736_  & \new_Sorter100|11737_ ;
  assign \new_Sorter100|11837_  = \new_Sorter100|11736_  | \new_Sorter100|11737_ ;
  assign \new_Sorter100|11838_  = \new_Sorter100|11738_  & \new_Sorter100|11739_ ;
  assign \new_Sorter100|11839_  = \new_Sorter100|11738_  | \new_Sorter100|11739_ ;
  assign \new_Sorter100|11840_  = \new_Sorter100|11740_  & \new_Sorter100|11741_ ;
  assign \new_Sorter100|11841_  = \new_Sorter100|11740_  | \new_Sorter100|11741_ ;
  assign \new_Sorter100|11842_  = \new_Sorter100|11742_  & \new_Sorter100|11743_ ;
  assign \new_Sorter100|11843_  = \new_Sorter100|11742_  | \new_Sorter100|11743_ ;
  assign \new_Sorter100|11844_  = \new_Sorter100|11744_  & \new_Sorter100|11745_ ;
  assign \new_Sorter100|11845_  = \new_Sorter100|11744_  | \new_Sorter100|11745_ ;
  assign \new_Sorter100|11846_  = \new_Sorter100|11746_  & \new_Sorter100|11747_ ;
  assign \new_Sorter100|11847_  = \new_Sorter100|11746_  | \new_Sorter100|11747_ ;
  assign \new_Sorter100|11848_  = \new_Sorter100|11748_  & \new_Sorter100|11749_ ;
  assign \new_Sorter100|11849_  = \new_Sorter100|11748_  | \new_Sorter100|11749_ ;
  assign \new_Sorter100|11850_  = \new_Sorter100|11750_  & \new_Sorter100|11751_ ;
  assign \new_Sorter100|11851_  = \new_Sorter100|11750_  | \new_Sorter100|11751_ ;
  assign \new_Sorter100|11852_  = \new_Sorter100|11752_  & \new_Sorter100|11753_ ;
  assign \new_Sorter100|11853_  = \new_Sorter100|11752_  | \new_Sorter100|11753_ ;
  assign \new_Sorter100|11854_  = \new_Sorter100|11754_  & \new_Sorter100|11755_ ;
  assign \new_Sorter100|11855_  = \new_Sorter100|11754_  | \new_Sorter100|11755_ ;
  assign \new_Sorter100|11856_  = \new_Sorter100|11756_  & \new_Sorter100|11757_ ;
  assign \new_Sorter100|11857_  = \new_Sorter100|11756_  | \new_Sorter100|11757_ ;
  assign \new_Sorter100|11858_  = \new_Sorter100|11758_  & \new_Sorter100|11759_ ;
  assign \new_Sorter100|11859_  = \new_Sorter100|11758_  | \new_Sorter100|11759_ ;
  assign \new_Sorter100|11860_  = \new_Sorter100|11760_  & \new_Sorter100|11761_ ;
  assign \new_Sorter100|11861_  = \new_Sorter100|11760_  | \new_Sorter100|11761_ ;
  assign \new_Sorter100|11862_  = \new_Sorter100|11762_  & \new_Sorter100|11763_ ;
  assign \new_Sorter100|11863_  = \new_Sorter100|11762_  | \new_Sorter100|11763_ ;
  assign \new_Sorter100|11864_  = \new_Sorter100|11764_  & \new_Sorter100|11765_ ;
  assign \new_Sorter100|11865_  = \new_Sorter100|11764_  | \new_Sorter100|11765_ ;
  assign \new_Sorter100|11866_  = \new_Sorter100|11766_  & \new_Sorter100|11767_ ;
  assign \new_Sorter100|11867_  = \new_Sorter100|11766_  | \new_Sorter100|11767_ ;
  assign \new_Sorter100|11868_  = \new_Sorter100|11768_  & \new_Sorter100|11769_ ;
  assign \new_Sorter100|11869_  = \new_Sorter100|11768_  | \new_Sorter100|11769_ ;
  assign \new_Sorter100|11870_  = \new_Sorter100|11770_  & \new_Sorter100|11771_ ;
  assign \new_Sorter100|11871_  = \new_Sorter100|11770_  | \new_Sorter100|11771_ ;
  assign \new_Sorter100|11872_  = \new_Sorter100|11772_  & \new_Sorter100|11773_ ;
  assign \new_Sorter100|11873_  = \new_Sorter100|11772_  | \new_Sorter100|11773_ ;
  assign \new_Sorter100|11874_  = \new_Sorter100|11774_  & \new_Sorter100|11775_ ;
  assign \new_Sorter100|11875_  = \new_Sorter100|11774_  | \new_Sorter100|11775_ ;
  assign \new_Sorter100|11876_  = \new_Sorter100|11776_  & \new_Sorter100|11777_ ;
  assign \new_Sorter100|11877_  = \new_Sorter100|11776_  | \new_Sorter100|11777_ ;
  assign \new_Sorter100|11878_  = \new_Sorter100|11778_  & \new_Sorter100|11779_ ;
  assign \new_Sorter100|11879_  = \new_Sorter100|11778_  | \new_Sorter100|11779_ ;
  assign \new_Sorter100|11880_  = \new_Sorter100|11780_  & \new_Sorter100|11781_ ;
  assign \new_Sorter100|11881_  = \new_Sorter100|11780_  | \new_Sorter100|11781_ ;
  assign \new_Sorter100|11882_  = \new_Sorter100|11782_  & \new_Sorter100|11783_ ;
  assign \new_Sorter100|11883_  = \new_Sorter100|11782_  | \new_Sorter100|11783_ ;
  assign \new_Sorter100|11884_  = \new_Sorter100|11784_  & \new_Sorter100|11785_ ;
  assign \new_Sorter100|11885_  = \new_Sorter100|11784_  | \new_Sorter100|11785_ ;
  assign \new_Sorter100|11886_  = \new_Sorter100|11786_  & \new_Sorter100|11787_ ;
  assign \new_Sorter100|11887_  = \new_Sorter100|11786_  | \new_Sorter100|11787_ ;
  assign \new_Sorter100|11888_  = \new_Sorter100|11788_  & \new_Sorter100|11789_ ;
  assign \new_Sorter100|11889_  = \new_Sorter100|11788_  | \new_Sorter100|11789_ ;
  assign \new_Sorter100|11890_  = \new_Sorter100|11790_  & \new_Sorter100|11791_ ;
  assign \new_Sorter100|11891_  = \new_Sorter100|11790_  | \new_Sorter100|11791_ ;
  assign \new_Sorter100|11892_  = \new_Sorter100|11792_  & \new_Sorter100|11793_ ;
  assign \new_Sorter100|11893_  = \new_Sorter100|11792_  | \new_Sorter100|11793_ ;
  assign \new_Sorter100|11894_  = \new_Sorter100|11794_  & \new_Sorter100|11795_ ;
  assign \new_Sorter100|11895_  = \new_Sorter100|11794_  | \new_Sorter100|11795_ ;
  assign \new_Sorter100|11896_  = \new_Sorter100|11796_  & \new_Sorter100|11797_ ;
  assign \new_Sorter100|11897_  = \new_Sorter100|11796_  | \new_Sorter100|11797_ ;
  assign \new_Sorter100|11898_  = \new_Sorter100|11798_  & \new_Sorter100|11799_ ;
  assign \new_Sorter100|11899_  = \new_Sorter100|11798_  | \new_Sorter100|11799_ ;
  assign \new_Sorter100|11900_  = \new_Sorter100|11800_ ;
  assign \new_Sorter100|11999_  = \new_Sorter100|11899_ ;
  assign \new_Sorter100|11901_  = \new_Sorter100|11801_  & \new_Sorter100|11802_ ;
  assign \new_Sorter100|11902_  = \new_Sorter100|11801_  | \new_Sorter100|11802_ ;
  assign \new_Sorter100|11903_  = \new_Sorter100|11803_  & \new_Sorter100|11804_ ;
  assign \new_Sorter100|11904_  = \new_Sorter100|11803_  | \new_Sorter100|11804_ ;
  assign \new_Sorter100|11905_  = \new_Sorter100|11805_  & \new_Sorter100|11806_ ;
  assign \new_Sorter100|11906_  = \new_Sorter100|11805_  | \new_Sorter100|11806_ ;
  assign \new_Sorter100|11907_  = \new_Sorter100|11807_  & \new_Sorter100|11808_ ;
  assign \new_Sorter100|11908_  = \new_Sorter100|11807_  | \new_Sorter100|11808_ ;
  assign \new_Sorter100|11909_  = \new_Sorter100|11809_  & \new_Sorter100|11810_ ;
  assign \new_Sorter100|11910_  = \new_Sorter100|11809_  | \new_Sorter100|11810_ ;
  assign \new_Sorter100|11911_  = \new_Sorter100|11811_  & \new_Sorter100|11812_ ;
  assign \new_Sorter100|11912_  = \new_Sorter100|11811_  | \new_Sorter100|11812_ ;
  assign \new_Sorter100|11913_  = \new_Sorter100|11813_  & \new_Sorter100|11814_ ;
  assign \new_Sorter100|11914_  = \new_Sorter100|11813_  | \new_Sorter100|11814_ ;
  assign \new_Sorter100|11915_  = \new_Sorter100|11815_  & \new_Sorter100|11816_ ;
  assign \new_Sorter100|11916_  = \new_Sorter100|11815_  | \new_Sorter100|11816_ ;
  assign \new_Sorter100|11917_  = \new_Sorter100|11817_  & \new_Sorter100|11818_ ;
  assign \new_Sorter100|11918_  = \new_Sorter100|11817_  | \new_Sorter100|11818_ ;
  assign \new_Sorter100|11919_  = \new_Sorter100|11819_  & \new_Sorter100|11820_ ;
  assign \new_Sorter100|11920_  = \new_Sorter100|11819_  | \new_Sorter100|11820_ ;
  assign \new_Sorter100|11921_  = \new_Sorter100|11821_  & \new_Sorter100|11822_ ;
  assign \new_Sorter100|11922_  = \new_Sorter100|11821_  | \new_Sorter100|11822_ ;
  assign \new_Sorter100|11923_  = \new_Sorter100|11823_  & \new_Sorter100|11824_ ;
  assign \new_Sorter100|11924_  = \new_Sorter100|11823_  | \new_Sorter100|11824_ ;
  assign \new_Sorter100|11925_  = \new_Sorter100|11825_  & \new_Sorter100|11826_ ;
  assign \new_Sorter100|11926_  = \new_Sorter100|11825_  | \new_Sorter100|11826_ ;
  assign \new_Sorter100|11927_  = \new_Sorter100|11827_  & \new_Sorter100|11828_ ;
  assign \new_Sorter100|11928_  = \new_Sorter100|11827_  | \new_Sorter100|11828_ ;
  assign \new_Sorter100|11929_  = \new_Sorter100|11829_  & \new_Sorter100|11830_ ;
  assign \new_Sorter100|11930_  = \new_Sorter100|11829_  | \new_Sorter100|11830_ ;
  assign \new_Sorter100|11931_  = \new_Sorter100|11831_  & \new_Sorter100|11832_ ;
  assign \new_Sorter100|11932_  = \new_Sorter100|11831_  | \new_Sorter100|11832_ ;
  assign \new_Sorter100|11933_  = \new_Sorter100|11833_  & \new_Sorter100|11834_ ;
  assign \new_Sorter100|11934_  = \new_Sorter100|11833_  | \new_Sorter100|11834_ ;
  assign \new_Sorter100|11935_  = \new_Sorter100|11835_  & \new_Sorter100|11836_ ;
  assign \new_Sorter100|11936_  = \new_Sorter100|11835_  | \new_Sorter100|11836_ ;
  assign \new_Sorter100|11937_  = \new_Sorter100|11837_  & \new_Sorter100|11838_ ;
  assign \new_Sorter100|11938_  = \new_Sorter100|11837_  | \new_Sorter100|11838_ ;
  assign \new_Sorter100|11939_  = \new_Sorter100|11839_  & \new_Sorter100|11840_ ;
  assign \new_Sorter100|11940_  = \new_Sorter100|11839_  | \new_Sorter100|11840_ ;
  assign \new_Sorter100|11941_  = \new_Sorter100|11841_  & \new_Sorter100|11842_ ;
  assign \new_Sorter100|11942_  = \new_Sorter100|11841_  | \new_Sorter100|11842_ ;
  assign \new_Sorter100|11943_  = \new_Sorter100|11843_  & \new_Sorter100|11844_ ;
  assign \new_Sorter100|11944_  = \new_Sorter100|11843_  | \new_Sorter100|11844_ ;
  assign \new_Sorter100|11945_  = \new_Sorter100|11845_  & \new_Sorter100|11846_ ;
  assign \new_Sorter100|11946_  = \new_Sorter100|11845_  | \new_Sorter100|11846_ ;
  assign \new_Sorter100|11947_  = \new_Sorter100|11847_  & \new_Sorter100|11848_ ;
  assign \new_Sorter100|11948_  = \new_Sorter100|11847_  | \new_Sorter100|11848_ ;
  assign \new_Sorter100|11949_  = \new_Sorter100|11849_  & \new_Sorter100|11850_ ;
  assign \new_Sorter100|11950_  = \new_Sorter100|11849_  | \new_Sorter100|11850_ ;
  assign \new_Sorter100|11951_  = \new_Sorter100|11851_  & \new_Sorter100|11852_ ;
  assign \new_Sorter100|11952_  = \new_Sorter100|11851_  | \new_Sorter100|11852_ ;
  assign \new_Sorter100|11953_  = \new_Sorter100|11853_  & \new_Sorter100|11854_ ;
  assign \new_Sorter100|11954_  = \new_Sorter100|11853_  | \new_Sorter100|11854_ ;
  assign \new_Sorter100|11955_  = \new_Sorter100|11855_  & \new_Sorter100|11856_ ;
  assign \new_Sorter100|11956_  = \new_Sorter100|11855_  | \new_Sorter100|11856_ ;
  assign \new_Sorter100|11957_  = \new_Sorter100|11857_  & \new_Sorter100|11858_ ;
  assign \new_Sorter100|11958_  = \new_Sorter100|11857_  | \new_Sorter100|11858_ ;
  assign \new_Sorter100|11959_  = \new_Sorter100|11859_  & \new_Sorter100|11860_ ;
  assign \new_Sorter100|11960_  = \new_Sorter100|11859_  | \new_Sorter100|11860_ ;
  assign \new_Sorter100|11961_  = \new_Sorter100|11861_  & \new_Sorter100|11862_ ;
  assign \new_Sorter100|11962_  = \new_Sorter100|11861_  | \new_Sorter100|11862_ ;
  assign \new_Sorter100|11963_  = \new_Sorter100|11863_  & \new_Sorter100|11864_ ;
  assign \new_Sorter100|11964_  = \new_Sorter100|11863_  | \new_Sorter100|11864_ ;
  assign \new_Sorter100|11965_  = \new_Sorter100|11865_  & \new_Sorter100|11866_ ;
  assign \new_Sorter100|11966_  = \new_Sorter100|11865_  | \new_Sorter100|11866_ ;
  assign \new_Sorter100|11967_  = \new_Sorter100|11867_  & \new_Sorter100|11868_ ;
  assign \new_Sorter100|11968_  = \new_Sorter100|11867_  | \new_Sorter100|11868_ ;
  assign \new_Sorter100|11969_  = \new_Sorter100|11869_  & \new_Sorter100|11870_ ;
  assign \new_Sorter100|11970_  = \new_Sorter100|11869_  | \new_Sorter100|11870_ ;
  assign \new_Sorter100|11971_  = \new_Sorter100|11871_  & \new_Sorter100|11872_ ;
  assign \new_Sorter100|11972_  = \new_Sorter100|11871_  | \new_Sorter100|11872_ ;
  assign \new_Sorter100|11973_  = \new_Sorter100|11873_  & \new_Sorter100|11874_ ;
  assign \new_Sorter100|11974_  = \new_Sorter100|11873_  | \new_Sorter100|11874_ ;
  assign \new_Sorter100|11975_  = \new_Sorter100|11875_  & \new_Sorter100|11876_ ;
  assign \new_Sorter100|11976_  = \new_Sorter100|11875_  | \new_Sorter100|11876_ ;
  assign \new_Sorter100|11977_  = \new_Sorter100|11877_  & \new_Sorter100|11878_ ;
  assign \new_Sorter100|11978_  = \new_Sorter100|11877_  | \new_Sorter100|11878_ ;
  assign \new_Sorter100|11979_  = \new_Sorter100|11879_  & \new_Sorter100|11880_ ;
  assign \new_Sorter100|11980_  = \new_Sorter100|11879_  | \new_Sorter100|11880_ ;
  assign \new_Sorter100|11981_  = \new_Sorter100|11881_  & \new_Sorter100|11882_ ;
  assign \new_Sorter100|11982_  = \new_Sorter100|11881_  | \new_Sorter100|11882_ ;
  assign \new_Sorter100|11983_  = \new_Sorter100|11883_  & \new_Sorter100|11884_ ;
  assign \new_Sorter100|11984_  = \new_Sorter100|11883_  | \new_Sorter100|11884_ ;
  assign \new_Sorter100|11985_  = \new_Sorter100|11885_  & \new_Sorter100|11886_ ;
  assign \new_Sorter100|11986_  = \new_Sorter100|11885_  | \new_Sorter100|11886_ ;
  assign \new_Sorter100|11987_  = \new_Sorter100|11887_  & \new_Sorter100|11888_ ;
  assign \new_Sorter100|11988_  = \new_Sorter100|11887_  | \new_Sorter100|11888_ ;
  assign \new_Sorter100|11989_  = \new_Sorter100|11889_  & \new_Sorter100|11890_ ;
  assign \new_Sorter100|11990_  = \new_Sorter100|11889_  | \new_Sorter100|11890_ ;
  assign \new_Sorter100|11991_  = \new_Sorter100|11891_  & \new_Sorter100|11892_ ;
  assign \new_Sorter100|11992_  = \new_Sorter100|11891_  | \new_Sorter100|11892_ ;
  assign \new_Sorter100|11993_  = \new_Sorter100|11893_  & \new_Sorter100|11894_ ;
  assign \new_Sorter100|11994_  = \new_Sorter100|11893_  | \new_Sorter100|11894_ ;
  assign \new_Sorter100|11995_  = \new_Sorter100|11895_  & \new_Sorter100|11896_ ;
  assign \new_Sorter100|11996_  = \new_Sorter100|11895_  | \new_Sorter100|11896_ ;
  assign \new_Sorter100|11997_  = \new_Sorter100|11897_  & \new_Sorter100|11898_ ;
  assign \new_Sorter100|11998_  = \new_Sorter100|11897_  | \new_Sorter100|11898_ ;
  assign \new_Sorter100|12000_  = \new_Sorter100|11900_  & \new_Sorter100|11901_ ;
  assign \new_Sorter100|12001_  = \new_Sorter100|11900_  | \new_Sorter100|11901_ ;
  assign \new_Sorter100|12002_  = \new_Sorter100|11902_  & \new_Sorter100|11903_ ;
  assign \new_Sorter100|12003_  = \new_Sorter100|11902_  | \new_Sorter100|11903_ ;
  assign \new_Sorter100|12004_  = \new_Sorter100|11904_  & \new_Sorter100|11905_ ;
  assign \new_Sorter100|12005_  = \new_Sorter100|11904_  | \new_Sorter100|11905_ ;
  assign \new_Sorter100|12006_  = \new_Sorter100|11906_  & \new_Sorter100|11907_ ;
  assign \new_Sorter100|12007_  = \new_Sorter100|11906_  | \new_Sorter100|11907_ ;
  assign \new_Sorter100|12008_  = \new_Sorter100|11908_  & \new_Sorter100|11909_ ;
  assign \new_Sorter100|12009_  = \new_Sorter100|11908_  | \new_Sorter100|11909_ ;
  assign \new_Sorter100|12010_  = \new_Sorter100|11910_  & \new_Sorter100|11911_ ;
  assign \new_Sorter100|12011_  = \new_Sorter100|11910_  | \new_Sorter100|11911_ ;
  assign \new_Sorter100|12012_  = \new_Sorter100|11912_  & \new_Sorter100|11913_ ;
  assign \new_Sorter100|12013_  = \new_Sorter100|11912_  | \new_Sorter100|11913_ ;
  assign \new_Sorter100|12014_  = \new_Sorter100|11914_  & \new_Sorter100|11915_ ;
  assign \new_Sorter100|12015_  = \new_Sorter100|11914_  | \new_Sorter100|11915_ ;
  assign \new_Sorter100|12016_  = \new_Sorter100|11916_  & \new_Sorter100|11917_ ;
  assign \new_Sorter100|12017_  = \new_Sorter100|11916_  | \new_Sorter100|11917_ ;
  assign \new_Sorter100|12018_  = \new_Sorter100|11918_  & \new_Sorter100|11919_ ;
  assign \new_Sorter100|12019_  = \new_Sorter100|11918_  | \new_Sorter100|11919_ ;
  assign \new_Sorter100|12020_  = \new_Sorter100|11920_  & \new_Sorter100|11921_ ;
  assign \new_Sorter100|12021_  = \new_Sorter100|11920_  | \new_Sorter100|11921_ ;
  assign \new_Sorter100|12022_  = \new_Sorter100|11922_  & \new_Sorter100|11923_ ;
  assign \new_Sorter100|12023_  = \new_Sorter100|11922_  | \new_Sorter100|11923_ ;
  assign \new_Sorter100|12024_  = \new_Sorter100|11924_  & \new_Sorter100|11925_ ;
  assign \new_Sorter100|12025_  = \new_Sorter100|11924_  | \new_Sorter100|11925_ ;
  assign \new_Sorter100|12026_  = \new_Sorter100|11926_  & \new_Sorter100|11927_ ;
  assign \new_Sorter100|12027_  = \new_Sorter100|11926_  | \new_Sorter100|11927_ ;
  assign \new_Sorter100|12028_  = \new_Sorter100|11928_  & \new_Sorter100|11929_ ;
  assign \new_Sorter100|12029_  = \new_Sorter100|11928_  | \new_Sorter100|11929_ ;
  assign \new_Sorter100|12030_  = \new_Sorter100|11930_  & \new_Sorter100|11931_ ;
  assign \new_Sorter100|12031_  = \new_Sorter100|11930_  | \new_Sorter100|11931_ ;
  assign \new_Sorter100|12032_  = \new_Sorter100|11932_  & \new_Sorter100|11933_ ;
  assign \new_Sorter100|12033_  = \new_Sorter100|11932_  | \new_Sorter100|11933_ ;
  assign \new_Sorter100|12034_  = \new_Sorter100|11934_  & \new_Sorter100|11935_ ;
  assign \new_Sorter100|12035_  = \new_Sorter100|11934_  | \new_Sorter100|11935_ ;
  assign \new_Sorter100|12036_  = \new_Sorter100|11936_  & \new_Sorter100|11937_ ;
  assign \new_Sorter100|12037_  = \new_Sorter100|11936_  | \new_Sorter100|11937_ ;
  assign \new_Sorter100|12038_  = \new_Sorter100|11938_  & \new_Sorter100|11939_ ;
  assign \new_Sorter100|12039_  = \new_Sorter100|11938_  | \new_Sorter100|11939_ ;
  assign \new_Sorter100|12040_  = \new_Sorter100|11940_  & \new_Sorter100|11941_ ;
  assign \new_Sorter100|12041_  = \new_Sorter100|11940_  | \new_Sorter100|11941_ ;
  assign \new_Sorter100|12042_  = \new_Sorter100|11942_  & \new_Sorter100|11943_ ;
  assign \new_Sorter100|12043_  = \new_Sorter100|11942_  | \new_Sorter100|11943_ ;
  assign \new_Sorter100|12044_  = \new_Sorter100|11944_  & \new_Sorter100|11945_ ;
  assign \new_Sorter100|12045_  = \new_Sorter100|11944_  | \new_Sorter100|11945_ ;
  assign \new_Sorter100|12046_  = \new_Sorter100|11946_  & \new_Sorter100|11947_ ;
  assign \new_Sorter100|12047_  = \new_Sorter100|11946_  | \new_Sorter100|11947_ ;
  assign \new_Sorter100|12048_  = \new_Sorter100|11948_  & \new_Sorter100|11949_ ;
  assign \new_Sorter100|12049_  = \new_Sorter100|11948_  | \new_Sorter100|11949_ ;
  assign \new_Sorter100|12050_  = \new_Sorter100|11950_  & \new_Sorter100|11951_ ;
  assign \new_Sorter100|12051_  = \new_Sorter100|11950_  | \new_Sorter100|11951_ ;
  assign \new_Sorter100|12052_  = \new_Sorter100|11952_  & \new_Sorter100|11953_ ;
  assign \new_Sorter100|12053_  = \new_Sorter100|11952_  | \new_Sorter100|11953_ ;
  assign \new_Sorter100|12054_  = \new_Sorter100|11954_  & \new_Sorter100|11955_ ;
  assign \new_Sorter100|12055_  = \new_Sorter100|11954_  | \new_Sorter100|11955_ ;
  assign \new_Sorter100|12056_  = \new_Sorter100|11956_  & \new_Sorter100|11957_ ;
  assign \new_Sorter100|12057_  = \new_Sorter100|11956_  | \new_Sorter100|11957_ ;
  assign \new_Sorter100|12058_  = \new_Sorter100|11958_  & \new_Sorter100|11959_ ;
  assign \new_Sorter100|12059_  = \new_Sorter100|11958_  | \new_Sorter100|11959_ ;
  assign \new_Sorter100|12060_  = \new_Sorter100|11960_  & \new_Sorter100|11961_ ;
  assign \new_Sorter100|12061_  = \new_Sorter100|11960_  | \new_Sorter100|11961_ ;
  assign \new_Sorter100|12062_  = \new_Sorter100|11962_  & \new_Sorter100|11963_ ;
  assign \new_Sorter100|12063_  = \new_Sorter100|11962_  | \new_Sorter100|11963_ ;
  assign \new_Sorter100|12064_  = \new_Sorter100|11964_  & \new_Sorter100|11965_ ;
  assign \new_Sorter100|12065_  = \new_Sorter100|11964_  | \new_Sorter100|11965_ ;
  assign \new_Sorter100|12066_  = \new_Sorter100|11966_  & \new_Sorter100|11967_ ;
  assign \new_Sorter100|12067_  = \new_Sorter100|11966_  | \new_Sorter100|11967_ ;
  assign \new_Sorter100|12068_  = \new_Sorter100|11968_  & \new_Sorter100|11969_ ;
  assign \new_Sorter100|12069_  = \new_Sorter100|11968_  | \new_Sorter100|11969_ ;
  assign \new_Sorter100|12070_  = \new_Sorter100|11970_  & \new_Sorter100|11971_ ;
  assign \new_Sorter100|12071_  = \new_Sorter100|11970_  | \new_Sorter100|11971_ ;
  assign \new_Sorter100|12072_  = \new_Sorter100|11972_  & \new_Sorter100|11973_ ;
  assign \new_Sorter100|12073_  = \new_Sorter100|11972_  | \new_Sorter100|11973_ ;
  assign \new_Sorter100|12074_  = \new_Sorter100|11974_  & \new_Sorter100|11975_ ;
  assign \new_Sorter100|12075_  = \new_Sorter100|11974_  | \new_Sorter100|11975_ ;
  assign \new_Sorter100|12076_  = \new_Sorter100|11976_  & \new_Sorter100|11977_ ;
  assign \new_Sorter100|12077_  = \new_Sorter100|11976_  | \new_Sorter100|11977_ ;
  assign \new_Sorter100|12078_  = \new_Sorter100|11978_  & \new_Sorter100|11979_ ;
  assign \new_Sorter100|12079_  = \new_Sorter100|11978_  | \new_Sorter100|11979_ ;
  assign \new_Sorter100|12080_  = \new_Sorter100|11980_  & \new_Sorter100|11981_ ;
  assign \new_Sorter100|12081_  = \new_Sorter100|11980_  | \new_Sorter100|11981_ ;
  assign \new_Sorter100|12082_  = \new_Sorter100|11982_  & \new_Sorter100|11983_ ;
  assign \new_Sorter100|12083_  = \new_Sorter100|11982_  | \new_Sorter100|11983_ ;
  assign \new_Sorter100|12084_  = \new_Sorter100|11984_  & \new_Sorter100|11985_ ;
  assign \new_Sorter100|12085_  = \new_Sorter100|11984_  | \new_Sorter100|11985_ ;
  assign \new_Sorter100|12086_  = \new_Sorter100|11986_  & \new_Sorter100|11987_ ;
  assign \new_Sorter100|12087_  = \new_Sorter100|11986_  | \new_Sorter100|11987_ ;
  assign \new_Sorter100|12088_  = \new_Sorter100|11988_  & \new_Sorter100|11989_ ;
  assign \new_Sorter100|12089_  = \new_Sorter100|11988_  | \new_Sorter100|11989_ ;
  assign \new_Sorter100|12090_  = \new_Sorter100|11990_  & \new_Sorter100|11991_ ;
  assign \new_Sorter100|12091_  = \new_Sorter100|11990_  | \new_Sorter100|11991_ ;
  assign \new_Sorter100|12092_  = \new_Sorter100|11992_  & \new_Sorter100|11993_ ;
  assign \new_Sorter100|12093_  = \new_Sorter100|11992_  | \new_Sorter100|11993_ ;
  assign \new_Sorter100|12094_  = \new_Sorter100|11994_  & \new_Sorter100|11995_ ;
  assign \new_Sorter100|12095_  = \new_Sorter100|11994_  | \new_Sorter100|11995_ ;
  assign \new_Sorter100|12096_  = \new_Sorter100|11996_  & \new_Sorter100|11997_ ;
  assign \new_Sorter100|12097_  = \new_Sorter100|11996_  | \new_Sorter100|11997_ ;
  assign \new_Sorter100|12098_  = \new_Sorter100|11998_  & \new_Sorter100|11999_ ;
  assign \new_Sorter100|12099_  = \new_Sorter100|11998_  | \new_Sorter100|11999_ ;
  assign \new_Sorter100|12100_  = \new_Sorter100|12000_ ;
  assign \new_Sorter100|12199_  = \new_Sorter100|12099_ ;
  assign \new_Sorter100|12101_  = \new_Sorter100|12001_  & \new_Sorter100|12002_ ;
  assign \new_Sorter100|12102_  = \new_Sorter100|12001_  | \new_Sorter100|12002_ ;
  assign \new_Sorter100|12103_  = \new_Sorter100|12003_  & \new_Sorter100|12004_ ;
  assign \new_Sorter100|12104_  = \new_Sorter100|12003_  | \new_Sorter100|12004_ ;
  assign \new_Sorter100|12105_  = \new_Sorter100|12005_  & \new_Sorter100|12006_ ;
  assign \new_Sorter100|12106_  = \new_Sorter100|12005_  | \new_Sorter100|12006_ ;
  assign \new_Sorter100|12107_  = \new_Sorter100|12007_  & \new_Sorter100|12008_ ;
  assign \new_Sorter100|12108_  = \new_Sorter100|12007_  | \new_Sorter100|12008_ ;
  assign \new_Sorter100|12109_  = \new_Sorter100|12009_  & \new_Sorter100|12010_ ;
  assign \new_Sorter100|12110_  = \new_Sorter100|12009_  | \new_Sorter100|12010_ ;
  assign \new_Sorter100|12111_  = \new_Sorter100|12011_  & \new_Sorter100|12012_ ;
  assign \new_Sorter100|12112_  = \new_Sorter100|12011_  | \new_Sorter100|12012_ ;
  assign \new_Sorter100|12113_  = \new_Sorter100|12013_  & \new_Sorter100|12014_ ;
  assign \new_Sorter100|12114_  = \new_Sorter100|12013_  | \new_Sorter100|12014_ ;
  assign \new_Sorter100|12115_  = \new_Sorter100|12015_  & \new_Sorter100|12016_ ;
  assign \new_Sorter100|12116_  = \new_Sorter100|12015_  | \new_Sorter100|12016_ ;
  assign \new_Sorter100|12117_  = \new_Sorter100|12017_  & \new_Sorter100|12018_ ;
  assign \new_Sorter100|12118_  = \new_Sorter100|12017_  | \new_Sorter100|12018_ ;
  assign \new_Sorter100|12119_  = \new_Sorter100|12019_  & \new_Sorter100|12020_ ;
  assign \new_Sorter100|12120_  = \new_Sorter100|12019_  | \new_Sorter100|12020_ ;
  assign \new_Sorter100|12121_  = \new_Sorter100|12021_  & \new_Sorter100|12022_ ;
  assign \new_Sorter100|12122_  = \new_Sorter100|12021_  | \new_Sorter100|12022_ ;
  assign \new_Sorter100|12123_  = \new_Sorter100|12023_  & \new_Sorter100|12024_ ;
  assign \new_Sorter100|12124_  = \new_Sorter100|12023_  | \new_Sorter100|12024_ ;
  assign \new_Sorter100|12125_  = \new_Sorter100|12025_  & \new_Sorter100|12026_ ;
  assign \new_Sorter100|12126_  = \new_Sorter100|12025_  | \new_Sorter100|12026_ ;
  assign \new_Sorter100|12127_  = \new_Sorter100|12027_  & \new_Sorter100|12028_ ;
  assign \new_Sorter100|12128_  = \new_Sorter100|12027_  | \new_Sorter100|12028_ ;
  assign \new_Sorter100|12129_  = \new_Sorter100|12029_  & \new_Sorter100|12030_ ;
  assign \new_Sorter100|12130_  = \new_Sorter100|12029_  | \new_Sorter100|12030_ ;
  assign \new_Sorter100|12131_  = \new_Sorter100|12031_  & \new_Sorter100|12032_ ;
  assign \new_Sorter100|12132_  = \new_Sorter100|12031_  | \new_Sorter100|12032_ ;
  assign \new_Sorter100|12133_  = \new_Sorter100|12033_  & \new_Sorter100|12034_ ;
  assign \new_Sorter100|12134_  = \new_Sorter100|12033_  | \new_Sorter100|12034_ ;
  assign \new_Sorter100|12135_  = \new_Sorter100|12035_  & \new_Sorter100|12036_ ;
  assign \new_Sorter100|12136_  = \new_Sorter100|12035_  | \new_Sorter100|12036_ ;
  assign \new_Sorter100|12137_  = \new_Sorter100|12037_  & \new_Sorter100|12038_ ;
  assign \new_Sorter100|12138_  = \new_Sorter100|12037_  | \new_Sorter100|12038_ ;
  assign \new_Sorter100|12139_  = \new_Sorter100|12039_  & \new_Sorter100|12040_ ;
  assign \new_Sorter100|12140_  = \new_Sorter100|12039_  | \new_Sorter100|12040_ ;
  assign \new_Sorter100|12141_  = \new_Sorter100|12041_  & \new_Sorter100|12042_ ;
  assign \new_Sorter100|12142_  = \new_Sorter100|12041_  | \new_Sorter100|12042_ ;
  assign \new_Sorter100|12143_  = \new_Sorter100|12043_  & \new_Sorter100|12044_ ;
  assign \new_Sorter100|12144_  = \new_Sorter100|12043_  | \new_Sorter100|12044_ ;
  assign \new_Sorter100|12145_  = \new_Sorter100|12045_  & \new_Sorter100|12046_ ;
  assign \new_Sorter100|12146_  = \new_Sorter100|12045_  | \new_Sorter100|12046_ ;
  assign \new_Sorter100|12147_  = \new_Sorter100|12047_  & \new_Sorter100|12048_ ;
  assign \new_Sorter100|12148_  = \new_Sorter100|12047_  | \new_Sorter100|12048_ ;
  assign \new_Sorter100|12149_  = \new_Sorter100|12049_  & \new_Sorter100|12050_ ;
  assign \new_Sorter100|12150_  = \new_Sorter100|12049_  | \new_Sorter100|12050_ ;
  assign \new_Sorter100|12151_  = \new_Sorter100|12051_  & \new_Sorter100|12052_ ;
  assign \new_Sorter100|12152_  = \new_Sorter100|12051_  | \new_Sorter100|12052_ ;
  assign \new_Sorter100|12153_  = \new_Sorter100|12053_  & \new_Sorter100|12054_ ;
  assign \new_Sorter100|12154_  = \new_Sorter100|12053_  | \new_Sorter100|12054_ ;
  assign \new_Sorter100|12155_  = \new_Sorter100|12055_  & \new_Sorter100|12056_ ;
  assign \new_Sorter100|12156_  = \new_Sorter100|12055_  | \new_Sorter100|12056_ ;
  assign \new_Sorter100|12157_  = \new_Sorter100|12057_  & \new_Sorter100|12058_ ;
  assign \new_Sorter100|12158_  = \new_Sorter100|12057_  | \new_Sorter100|12058_ ;
  assign \new_Sorter100|12159_  = \new_Sorter100|12059_  & \new_Sorter100|12060_ ;
  assign \new_Sorter100|12160_  = \new_Sorter100|12059_  | \new_Sorter100|12060_ ;
  assign \new_Sorter100|12161_  = \new_Sorter100|12061_  & \new_Sorter100|12062_ ;
  assign \new_Sorter100|12162_  = \new_Sorter100|12061_  | \new_Sorter100|12062_ ;
  assign \new_Sorter100|12163_  = \new_Sorter100|12063_  & \new_Sorter100|12064_ ;
  assign \new_Sorter100|12164_  = \new_Sorter100|12063_  | \new_Sorter100|12064_ ;
  assign \new_Sorter100|12165_  = \new_Sorter100|12065_  & \new_Sorter100|12066_ ;
  assign \new_Sorter100|12166_  = \new_Sorter100|12065_  | \new_Sorter100|12066_ ;
  assign \new_Sorter100|12167_  = \new_Sorter100|12067_  & \new_Sorter100|12068_ ;
  assign \new_Sorter100|12168_  = \new_Sorter100|12067_  | \new_Sorter100|12068_ ;
  assign \new_Sorter100|12169_  = \new_Sorter100|12069_  & \new_Sorter100|12070_ ;
  assign \new_Sorter100|12170_  = \new_Sorter100|12069_  | \new_Sorter100|12070_ ;
  assign \new_Sorter100|12171_  = \new_Sorter100|12071_  & \new_Sorter100|12072_ ;
  assign \new_Sorter100|12172_  = \new_Sorter100|12071_  | \new_Sorter100|12072_ ;
  assign \new_Sorter100|12173_  = \new_Sorter100|12073_  & \new_Sorter100|12074_ ;
  assign \new_Sorter100|12174_  = \new_Sorter100|12073_  | \new_Sorter100|12074_ ;
  assign \new_Sorter100|12175_  = \new_Sorter100|12075_  & \new_Sorter100|12076_ ;
  assign \new_Sorter100|12176_  = \new_Sorter100|12075_  | \new_Sorter100|12076_ ;
  assign \new_Sorter100|12177_  = \new_Sorter100|12077_  & \new_Sorter100|12078_ ;
  assign \new_Sorter100|12178_  = \new_Sorter100|12077_  | \new_Sorter100|12078_ ;
  assign \new_Sorter100|12179_  = \new_Sorter100|12079_  & \new_Sorter100|12080_ ;
  assign \new_Sorter100|12180_  = \new_Sorter100|12079_  | \new_Sorter100|12080_ ;
  assign \new_Sorter100|12181_  = \new_Sorter100|12081_  & \new_Sorter100|12082_ ;
  assign \new_Sorter100|12182_  = \new_Sorter100|12081_  | \new_Sorter100|12082_ ;
  assign \new_Sorter100|12183_  = \new_Sorter100|12083_  & \new_Sorter100|12084_ ;
  assign \new_Sorter100|12184_  = \new_Sorter100|12083_  | \new_Sorter100|12084_ ;
  assign \new_Sorter100|12185_  = \new_Sorter100|12085_  & \new_Sorter100|12086_ ;
  assign \new_Sorter100|12186_  = \new_Sorter100|12085_  | \new_Sorter100|12086_ ;
  assign \new_Sorter100|12187_  = \new_Sorter100|12087_  & \new_Sorter100|12088_ ;
  assign \new_Sorter100|12188_  = \new_Sorter100|12087_  | \new_Sorter100|12088_ ;
  assign \new_Sorter100|12189_  = \new_Sorter100|12089_  & \new_Sorter100|12090_ ;
  assign \new_Sorter100|12190_  = \new_Sorter100|12089_  | \new_Sorter100|12090_ ;
  assign \new_Sorter100|12191_  = \new_Sorter100|12091_  & \new_Sorter100|12092_ ;
  assign \new_Sorter100|12192_  = \new_Sorter100|12091_  | \new_Sorter100|12092_ ;
  assign \new_Sorter100|12193_  = \new_Sorter100|12093_  & \new_Sorter100|12094_ ;
  assign \new_Sorter100|12194_  = \new_Sorter100|12093_  | \new_Sorter100|12094_ ;
  assign \new_Sorter100|12195_  = \new_Sorter100|12095_  & \new_Sorter100|12096_ ;
  assign \new_Sorter100|12196_  = \new_Sorter100|12095_  | \new_Sorter100|12096_ ;
  assign \new_Sorter100|12197_  = \new_Sorter100|12097_  & \new_Sorter100|12098_ ;
  assign \new_Sorter100|12198_  = \new_Sorter100|12097_  | \new_Sorter100|12098_ ;
  assign \new_Sorter100|12200_  = \new_Sorter100|12100_  & \new_Sorter100|12101_ ;
  assign \new_Sorter100|12201_  = \new_Sorter100|12100_  | \new_Sorter100|12101_ ;
  assign \new_Sorter100|12202_  = \new_Sorter100|12102_  & \new_Sorter100|12103_ ;
  assign \new_Sorter100|12203_  = \new_Sorter100|12102_  | \new_Sorter100|12103_ ;
  assign \new_Sorter100|12204_  = \new_Sorter100|12104_  & \new_Sorter100|12105_ ;
  assign \new_Sorter100|12205_  = \new_Sorter100|12104_  | \new_Sorter100|12105_ ;
  assign \new_Sorter100|12206_  = \new_Sorter100|12106_  & \new_Sorter100|12107_ ;
  assign \new_Sorter100|12207_  = \new_Sorter100|12106_  | \new_Sorter100|12107_ ;
  assign \new_Sorter100|12208_  = \new_Sorter100|12108_  & \new_Sorter100|12109_ ;
  assign \new_Sorter100|12209_  = \new_Sorter100|12108_  | \new_Sorter100|12109_ ;
  assign \new_Sorter100|12210_  = \new_Sorter100|12110_  & \new_Sorter100|12111_ ;
  assign \new_Sorter100|12211_  = \new_Sorter100|12110_  | \new_Sorter100|12111_ ;
  assign \new_Sorter100|12212_  = \new_Sorter100|12112_  & \new_Sorter100|12113_ ;
  assign \new_Sorter100|12213_  = \new_Sorter100|12112_  | \new_Sorter100|12113_ ;
  assign \new_Sorter100|12214_  = \new_Sorter100|12114_  & \new_Sorter100|12115_ ;
  assign \new_Sorter100|12215_  = \new_Sorter100|12114_  | \new_Sorter100|12115_ ;
  assign \new_Sorter100|12216_  = \new_Sorter100|12116_  & \new_Sorter100|12117_ ;
  assign \new_Sorter100|12217_  = \new_Sorter100|12116_  | \new_Sorter100|12117_ ;
  assign \new_Sorter100|12218_  = \new_Sorter100|12118_  & \new_Sorter100|12119_ ;
  assign \new_Sorter100|12219_  = \new_Sorter100|12118_  | \new_Sorter100|12119_ ;
  assign \new_Sorter100|12220_  = \new_Sorter100|12120_  & \new_Sorter100|12121_ ;
  assign \new_Sorter100|12221_  = \new_Sorter100|12120_  | \new_Sorter100|12121_ ;
  assign \new_Sorter100|12222_  = \new_Sorter100|12122_  & \new_Sorter100|12123_ ;
  assign \new_Sorter100|12223_  = \new_Sorter100|12122_  | \new_Sorter100|12123_ ;
  assign \new_Sorter100|12224_  = \new_Sorter100|12124_  & \new_Sorter100|12125_ ;
  assign \new_Sorter100|12225_  = \new_Sorter100|12124_  | \new_Sorter100|12125_ ;
  assign \new_Sorter100|12226_  = \new_Sorter100|12126_  & \new_Sorter100|12127_ ;
  assign \new_Sorter100|12227_  = \new_Sorter100|12126_  | \new_Sorter100|12127_ ;
  assign \new_Sorter100|12228_  = \new_Sorter100|12128_  & \new_Sorter100|12129_ ;
  assign \new_Sorter100|12229_  = \new_Sorter100|12128_  | \new_Sorter100|12129_ ;
  assign \new_Sorter100|12230_  = \new_Sorter100|12130_  & \new_Sorter100|12131_ ;
  assign \new_Sorter100|12231_  = \new_Sorter100|12130_  | \new_Sorter100|12131_ ;
  assign \new_Sorter100|12232_  = \new_Sorter100|12132_  & \new_Sorter100|12133_ ;
  assign \new_Sorter100|12233_  = \new_Sorter100|12132_  | \new_Sorter100|12133_ ;
  assign \new_Sorter100|12234_  = \new_Sorter100|12134_  & \new_Sorter100|12135_ ;
  assign \new_Sorter100|12235_  = \new_Sorter100|12134_  | \new_Sorter100|12135_ ;
  assign \new_Sorter100|12236_  = \new_Sorter100|12136_  & \new_Sorter100|12137_ ;
  assign \new_Sorter100|12237_  = \new_Sorter100|12136_  | \new_Sorter100|12137_ ;
  assign \new_Sorter100|12238_  = \new_Sorter100|12138_  & \new_Sorter100|12139_ ;
  assign \new_Sorter100|12239_  = \new_Sorter100|12138_  | \new_Sorter100|12139_ ;
  assign \new_Sorter100|12240_  = \new_Sorter100|12140_  & \new_Sorter100|12141_ ;
  assign \new_Sorter100|12241_  = \new_Sorter100|12140_  | \new_Sorter100|12141_ ;
  assign \new_Sorter100|12242_  = \new_Sorter100|12142_  & \new_Sorter100|12143_ ;
  assign \new_Sorter100|12243_  = \new_Sorter100|12142_  | \new_Sorter100|12143_ ;
  assign \new_Sorter100|12244_  = \new_Sorter100|12144_  & \new_Sorter100|12145_ ;
  assign \new_Sorter100|12245_  = \new_Sorter100|12144_  | \new_Sorter100|12145_ ;
  assign \new_Sorter100|12246_  = \new_Sorter100|12146_  & \new_Sorter100|12147_ ;
  assign \new_Sorter100|12247_  = \new_Sorter100|12146_  | \new_Sorter100|12147_ ;
  assign \new_Sorter100|12248_  = \new_Sorter100|12148_  & \new_Sorter100|12149_ ;
  assign \new_Sorter100|12249_  = \new_Sorter100|12148_  | \new_Sorter100|12149_ ;
  assign \new_Sorter100|12250_  = \new_Sorter100|12150_  & \new_Sorter100|12151_ ;
  assign \new_Sorter100|12251_  = \new_Sorter100|12150_  | \new_Sorter100|12151_ ;
  assign \new_Sorter100|12252_  = \new_Sorter100|12152_  & \new_Sorter100|12153_ ;
  assign \new_Sorter100|12253_  = \new_Sorter100|12152_  | \new_Sorter100|12153_ ;
  assign \new_Sorter100|12254_  = \new_Sorter100|12154_  & \new_Sorter100|12155_ ;
  assign \new_Sorter100|12255_  = \new_Sorter100|12154_  | \new_Sorter100|12155_ ;
  assign \new_Sorter100|12256_  = \new_Sorter100|12156_  & \new_Sorter100|12157_ ;
  assign \new_Sorter100|12257_  = \new_Sorter100|12156_  | \new_Sorter100|12157_ ;
  assign \new_Sorter100|12258_  = \new_Sorter100|12158_  & \new_Sorter100|12159_ ;
  assign \new_Sorter100|12259_  = \new_Sorter100|12158_  | \new_Sorter100|12159_ ;
  assign \new_Sorter100|12260_  = \new_Sorter100|12160_  & \new_Sorter100|12161_ ;
  assign \new_Sorter100|12261_  = \new_Sorter100|12160_  | \new_Sorter100|12161_ ;
  assign \new_Sorter100|12262_  = \new_Sorter100|12162_  & \new_Sorter100|12163_ ;
  assign \new_Sorter100|12263_  = \new_Sorter100|12162_  | \new_Sorter100|12163_ ;
  assign \new_Sorter100|12264_  = \new_Sorter100|12164_  & \new_Sorter100|12165_ ;
  assign \new_Sorter100|12265_  = \new_Sorter100|12164_  | \new_Sorter100|12165_ ;
  assign \new_Sorter100|12266_  = \new_Sorter100|12166_  & \new_Sorter100|12167_ ;
  assign \new_Sorter100|12267_  = \new_Sorter100|12166_  | \new_Sorter100|12167_ ;
  assign \new_Sorter100|12268_  = \new_Sorter100|12168_  & \new_Sorter100|12169_ ;
  assign \new_Sorter100|12269_  = \new_Sorter100|12168_  | \new_Sorter100|12169_ ;
  assign \new_Sorter100|12270_  = \new_Sorter100|12170_  & \new_Sorter100|12171_ ;
  assign \new_Sorter100|12271_  = \new_Sorter100|12170_  | \new_Sorter100|12171_ ;
  assign \new_Sorter100|12272_  = \new_Sorter100|12172_  & \new_Sorter100|12173_ ;
  assign \new_Sorter100|12273_  = \new_Sorter100|12172_  | \new_Sorter100|12173_ ;
  assign \new_Sorter100|12274_  = \new_Sorter100|12174_  & \new_Sorter100|12175_ ;
  assign \new_Sorter100|12275_  = \new_Sorter100|12174_  | \new_Sorter100|12175_ ;
  assign \new_Sorter100|12276_  = \new_Sorter100|12176_  & \new_Sorter100|12177_ ;
  assign \new_Sorter100|12277_  = \new_Sorter100|12176_  | \new_Sorter100|12177_ ;
  assign \new_Sorter100|12278_  = \new_Sorter100|12178_  & \new_Sorter100|12179_ ;
  assign \new_Sorter100|12279_  = \new_Sorter100|12178_  | \new_Sorter100|12179_ ;
  assign \new_Sorter100|12280_  = \new_Sorter100|12180_  & \new_Sorter100|12181_ ;
  assign \new_Sorter100|12281_  = \new_Sorter100|12180_  | \new_Sorter100|12181_ ;
  assign \new_Sorter100|12282_  = \new_Sorter100|12182_  & \new_Sorter100|12183_ ;
  assign \new_Sorter100|12283_  = \new_Sorter100|12182_  | \new_Sorter100|12183_ ;
  assign \new_Sorter100|12284_  = \new_Sorter100|12184_  & \new_Sorter100|12185_ ;
  assign \new_Sorter100|12285_  = \new_Sorter100|12184_  | \new_Sorter100|12185_ ;
  assign \new_Sorter100|12286_  = \new_Sorter100|12186_  & \new_Sorter100|12187_ ;
  assign \new_Sorter100|12287_  = \new_Sorter100|12186_  | \new_Sorter100|12187_ ;
  assign \new_Sorter100|12288_  = \new_Sorter100|12188_  & \new_Sorter100|12189_ ;
  assign \new_Sorter100|12289_  = \new_Sorter100|12188_  | \new_Sorter100|12189_ ;
  assign \new_Sorter100|12290_  = \new_Sorter100|12190_  & \new_Sorter100|12191_ ;
  assign \new_Sorter100|12291_  = \new_Sorter100|12190_  | \new_Sorter100|12191_ ;
  assign \new_Sorter100|12292_  = \new_Sorter100|12192_  & \new_Sorter100|12193_ ;
  assign \new_Sorter100|12293_  = \new_Sorter100|12192_  | \new_Sorter100|12193_ ;
  assign \new_Sorter100|12294_  = \new_Sorter100|12194_  & \new_Sorter100|12195_ ;
  assign \new_Sorter100|12295_  = \new_Sorter100|12194_  | \new_Sorter100|12195_ ;
  assign \new_Sorter100|12296_  = \new_Sorter100|12196_  & \new_Sorter100|12197_ ;
  assign \new_Sorter100|12297_  = \new_Sorter100|12196_  | \new_Sorter100|12197_ ;
  assign \new_Sorter100|12298_  = \new_Sorter100|12198_  & \new_Sorter100|12199_ ;
  assign \new_Sorter100|12299_  = \new_Sorter100|12198_  | \new_Sorter100|12199_ ;
  assign \new_Sorter100|12300_  = \new_Sorter100|12200_ ;
  assign \new_Sorter100|12399_  = \new_Sorter100|12299_ ;
  assign \new_Sorter100|12301_  = \new_Sorter100|12201_  & \new_Sorter100|12202_ ;
  assign \new_Sorter100|12302_  = \new_Sorter100|12201_  | \new_Sorter100|12202_ ;
  assign \new_Sorter100|12303_  = \new_Sorter100|12203_  & \new_Sorter100|12204_ ;
  assign \new_Sorter100|12304_  = \new_Sorter100|12203_  | \new_Sorter100|12204_ ;
  assign \new_Sorter100|12305_  = \new_Sorter100|12205_  & \new_Sorter100|12206_ ;
  assign \new_Sorter100|12306_  = \new_Sorter100|12205_  | \new_Sorter100|12206_ ;
  assign \new_Sorter100|12307_  = \new_Sorter100|12207_  & \new_Sorter100|12208_ ;
  assign \new_Sorter100|12308_  = \new_Sorter100|12207_  | \new_Sorter100|12208_ ;
  assign \new_Sorter100|12309_  = \new_Sorter100|12209_  & \new_Sorter100|12210_ ;
  assign \new_Sorter100|12310_  = \new_Sorter100|12209_  | \new_Sorter100|12210_ ;
  assign \new_Sorter100|12311_  = \new_Sorter100|12211_  & \new_Sorter100|12212_ ;
  assign \new_Sorter100|12312_  = \new_Sorter100|12211_  | \new_Sorter100|12212_ ;
  assign \new_Sorter100|12313_  = \new_Sorter100|12213_  & \new_Sorter100|12214_ ;
  assign \new_Sorter100|12314_  = \new_Sorter100|12213_  | \new_Sorter100|12214_ ;
  assign \new_Sorter100|12315_  = \new_Sorter100|12215_  & \new_Sorter100|12216_ ;
  assign \new_Sorter100|12316_  = \new_Sorter100|12215_  | \new_Sorter100|12216_ ;
  assign \new_Sorter100|12317_  = \new_Sorter100|12217_  & \new_Sorter100|12218_ ;
  assign \new_Sorter100|12318_  = \new_Sorter100|12217_  | \new_Sorter100|12218_ ;
  assign \new_Sorter100|12319_  = \new_Sorter100|12219_  & \new_Sorter100|12220_ ;
  assign \new_Sorter100|12320_  = \new_Sorter100|12219_  | \new_Sorter100|12220_ ;
  assign \new_Sorter100|12321_  = \new_Sorter100|12221_  & \new_Sorter100|12222_ ;
  assign \new_Sorter100|12322_  = \new_Sorter100|12221_  | \new_Sorter100|12222_ ;
  assign \new_Sorter100|12323_  = \new_Sorter100|12223_  & \new_Sorter100|12224_ ;
  assign \new_Sorter100|12324_  = \new_Sorter100|12223_  | \new_Sorter100|12224_ ;
  assign \new_Sorter100|12325_  = \new_Sorter100|12225_  & \new_Sorter100|12226_ ;
  assign \new_Sorter100|12326_  = \new_Sorter100|12225_  | \new_Sorter100|12226_ ;
  assign \new_Sorter100|12327_  = \new_Sorter100|12227_  & \new_Sorter100|12228_ ;
  assign \new_Sorter100|12328_  = \new_Sorter100|12227_  | \new_Sorter100|12228_ ;
  assign \new_Sorter100|12329_  = \new_Sorter100|12229_  & \new_Sorter100|12230_ ;
  assign \new_Sorter100|12330_  = \new_Sorter100|12229_  | \new_Sorter100|12230_ ;
  assign \new_Sorter100|12331_  = \new_Sorter100|12231_  & \new_Sorter100|12232_ ;
  assign \new_Sorter100|12332_  = \new_Sorter100|12231_  | \new_Sorter100|12232_ ;
  assign \new_Sorter100|12333_  = \new_Sorter100|12233_  & \new_Sorter100|12234_ ;
  assign \new_Sorter100|12334_  = \new_Sorter100|12233_  | \new_Sorter100|12234_ ;
  assign \new_Sorter100|12335_  = \new_Sorter100|12235_  & \new_Sorter100|12236_ ;
  assign \new_Sorter100|12336_  = \new_Sorter100|12235_  | \new_Sorter100|12236_ ;
  assign \new_Sorter100|12337_  = \new_Sorter100|12237_  & \new_Sorter100|12238_ ;
  assign \new_Sorter100|12338_  = \new_Sorter100|12237_  | \new_Sorter100|12238_ ;
  assign \new_Sorter100|12339_  = \new_Sorter100|12239_  & \new_Sorter100|12240_ ;
  assign \new_Sorter100|12340_  = \new_Sorter100|12239_  | \new_Sorter100|12240_ ;
  assign \new_Sorter100|12341_  = \new_Sorter100|12241_  & \new_Sorter100|12242_ ;
  assign \new_Sorter100|12342_  = \new_Sorter100|12241_  | \new_Sorter100|12242_ ;
  assign \new_Sorter100|12343_  = \new_Sorter100|12243_  & \new_Sorter100|12244_ ;
  assign \new_Sorter100|12344_  = \new_Sorter100|12243_  | \new_Sorter100|12244_ ;
  assign \new_Sorter100|12345_  = \new_Sorter100|12245_  & \new_Sorter100|12246_ ;
  assign \new_Sorter100|12346_  = \new_Sorter100|12245_  | \new_Sorter100|12246_ ;
  assign \new_Sorter100|12347_  = \new_Sorter100|12247_  & \new_Sorter100|12248_ ;
  assign \new_Sorter100|12348_  = \new_Sorter100|12247_  | \new_Sorter100|12248_ ;
  assign \new_Sorter100|12349_  = \new_Sorter100|12249_  & \new_Sorter100|12250_ ;
  assign \new_Sorter100|12350_  = \new_Sorter100|12249_  | \new_Sorter100|12250_ ;
  assign \new_Sorter100|12351_  = \new_Sorter100|12251_  & \new_Sorter100|12252_ ;
  assign \new_Sorter100|12352_  = \new_Sorter100|12251_  | \new_Sorter100|12252_ ;
  assign \new_Sorter100|12353_  = \new_Sorter100|12253_  & \new_Sorter100|12254_ ;
  assign \new_Sorter100|12354_  = \new_Sorter100|12253_  | \new_Sorter100|12254_ ;
  assign \new_Sorter100|12355_  = \new_Sorter100|12255_  & \new_Sorter100|12256_ ;
  assign \new_Sorter100|12356_  = \new_Sorter100|12255_  | \new_Sorter100|12256_ ;
  assign \new_Sorter100|12357_  = \new_Sorter100|12257_  & \new_Sorter100|12258_ ;
  assign \new_Sorter100|12358_  = \new_Sorter100|12257_  | \new_Sorter100|12258_ ;
  assign \new_Sorter100|12359_  = \new_Sorter100|12259_  & \new_Sorter100|12260_ ;
  assign \new_Sorter100|12360_  = \new_Sorter100|12259_  | \new_Sorter100|12260_ ;
  assign \new_Sorter100|12361_  = \new_Sorter100|12261_  & \new_Sorter100|12262_ ;
  assign \new_Sorter100|12362_  = \new_Sorter100|12261_  | \new_Sorter100|12262_ ;
  assign \new_Sorter100|12363_  = \new_Sorter100|12263_  & \new_Sorter100|12264_ ;
  assign \new_Sorter100|12364_  = \new_Sorter100|12263_  | \new_Sorter100|12264_ ;
  assign \new_Sorter100|12365_  = \new_Sorter100|12265_  & \new_Sorter100|12266_ ;
  assign \new_Sorter100|12366_  = \new_Sorter100|12265_  | \new_Sorter100|12266_ ;
  assign \new_Sorter100|12367_  = \new_Sorter100|12267_  & \new_Sorter100|12268_ ;
  assign \new_Sorter100|12368_  = \new_Sorter100|12267_  | \new_Sorter100|12268_ ;
  assign \new_Sorter100|12369_  = \new_Sorter100|12269_  & \new_Sorter100|12270_ ;
  assign \new_Sorter100|12370_  = \new_Sorter100|12269_  | \new_Sorter100|12270_ ;
  assign \new_Sorter100|12371_  = \new_Sorter100|12271_  & \new_Sorter100|12272_ ;
  assign \new_Sorter100|12372_  = \new_Sorter100|12271_  | \new_Sorter100|12272_ ;
  assign \new_Sorter100|12373_  = \new_Sorter100|12273_  & \new_Sorter100|12274_ ;
  assign \new_Sorter100|12374_  = \new_Sorter100|12273_  | \new_Sorter100|12274_ ;
  assign \new_Sorter100|12375_  = \new_Sorter100|12275_  & \new_Sorter100|12276_ ;
  assign \new_Sorter100|12376_  = \new_Sorter100|12275_  | \new_Sorter100|12276_ ;
  assign \new_Sorter100|12377_  = \new_Sorter100|12277_  & \new_Sorter100|12278_ ;
  assign \new_Sorter100|12378_  = \new_Sorter100|12277_  | \new_Sorter100|12278_ ;
  assign \new_Sorter100|12379_  = \new_Sorter100|12279_  & \new_Sorter100|12280_ ;
  assign \new_Sorter100|12380_  = \new_Sorter100|12279_  | \new_Sorter100|12280_ ;
  assign \new_Sorter100|12381_  = \new_Sorter100|12281_  & \new_Sorter100|12282_ ;
  assign \new_Sorter100|12382_  = \new_Sorter100|12281_  | \new_Sorter100|12282_ ;
  assign \new_Sorter100|12383_  = \new_Sorter100|12283_  & \new_Sorter100|12284_ ;
  assign \new_Sorter100|12384_  = \new_Sorter100|12283_  | \new_Sorter100|12284_ ;
  assign \new_Sorter100|12385_  = \new_Sorter100|12285_  & \new_Sorter100|12286_ ;
  assign \new_Sorter100|12386_  = \new_Sorter100|12285_  | \new_Sorter100|12286_ ;
  assign \new_Sorter100|12387_  = \new_Sorter100|12287_  & \new_Sorter100|12288_ ;
  assign \new_Sorter100|12388_  = \new_Sorter100|12287_  | \new_Sorter100|12288_ ;
  assign \new_Sorter100|12389_  = \new_Sorter100|12289_  & \new_Sorter100|12290_ ;
  assign \new_Sorter100|12390_  = \new_Sorter100|12289_  | \new_Sorter100|12290_ ;
  assign \new_Sorter100|12391_  = \new_Sorter100|12291_  & \new_Sorter100|12292_ ;
  assign \new_Sorter100|12392_  = \new_Sorter100|12291_  | \new_Sorter100|12292_ ;
  assign \new_Sorter100|12393_  = \new_Sorter100|12293_  & \new_Sorter100|12294_ ;
  assign \new_Sorter100|12394_  = \new_Sorter100|12293_  | \new_Sorter100|12294_ ;
  assign \new_Sorter100|12395_  = \new_Sorter100|12295_  & \new_Sorter100|12296_ ;
  assign \new_Sorter100|12396_  = \new_Sorter100|12295_  | \new_Sorter100|12296_ ;
  assign \new_Sorter100|12397_  = \new_Sorter100|12297_  & \new_Sorter100|12298_ ;
  assign \new_Sorter100|12398_  = \new_Sorter100|12297_  | \new_Sorter100|12298_ ;
  assign \new_Sorter100|12400_  = \new_Sorter100|12300_  & \new_Sorter100|12301_ ;
  assign \new_Sorter100|12401_  = \new_Sorter100|12300_  | \new_Sorter100|12301_ ;
  assign \new_Sorter100|12402_  = \new_Sorter100|12302_  & \new_Sorter100|12303_ ;
  assign \new_Sorter100|12403_  = \new_Sorter100|12302_  | \new_Sorter100|12303_ ;
  assign \new_Sorter100|12404_  = \new_Sorter100|12304_  & \new_Sorter100|12305_ ;
  assign \new_Sorter100|12405_  = \new_Sorter100|12304_  | \new_Sorter100|12305_ ;
  assign \new_Sorter100|12406_  = \new_Sorter100|12306_  & \new_Sorter100|12307_ ;
  assign \new_Sorter100|12407_  = \new_Sorter100|12306_  | \new_Sorter100|12307_ ;
  assign \new_Sorter100|12408_  = \new_Sorter100|12308_  & \new_Sorter100|12309_ ;
  assign \new_Sorter100|12409_  = \new_Sorter100|12308_  | \new_Sorter100|12309_ ;
  assign \new_Sorter100|12410_  = \new_Sorter100|12310_  & \new_Sorter100|12311_ ;
  assign \new_Sorter100|12411_  = \new_Sorter100|12310_  | \new_Sorter100|12311_ ;
  assign \new_Sorter100|12412_  = \new_Sorter100|12312_  & \new_Sorter100|12313_ ;
  assign \new_Sorter100|12413_  = \new_Sorter100|12312_  | \new_Sorter100|12313_ ;
  assign \new_Sorter100|12414_  = \new_Sorter100|12314_  & \new_Sorter100|12315_ ;
  assign \new_Sorter100|12415_  = \new_Sorter100|12314_  | \new_Sorter100|12315_ ;
  assign \new_Sorter100|12416_  = \new_Sorter100|12316_  & \new_Sorter100|12317_ ;
  assign \new_Sorter100|12417_  = \new_Sorter100|12316_  | \new_Sorter100|12317_ ;
  assign \new_Sorter100|12418_  = \new_Sorter100|12318_  & \new_Sorter100|12319_ ;
  assign \new_Sorter100|12419_  = \new_Sorter100|12318_  | \new_Sorter100|12319_ ;
  assign \new_Sorter100|12420_  = \new_Sorter100|12320_  & \new_Sorter100|12321_ ;
  assign \new_Sorter100|12421_  = \new_Sorter100|12320_  | \new_Sorter100|12321_ ;
  assign \new_Sorter100|12422_  = \new_Sorter100|12322_  & \new_Sorter100|12323_ ;
  assign \new_Sorter100|12423_  = \new_Sorter100|12322_  | \new_Sorter100|12323_ ;
  assign \new_Sorter100|12424_  = \new_Sorter100|12324_  & \new_Sorter100|12325_ ;
  assign \new_Sorter100|12425_  = \new_Sorter100|12324_  | \new_Sorter100|12325_ ;
  assign \new_Sorter100|12426_  = \new_Sorter100|12326_  & \new_Sorter100|12327_ ;
  assign \new_Sorter100|12427_  = \new_Sorter100|12326_  | \new_Sorter100|12327_ ;
  assign \new_Sorter100|12428_  = \new_Sorter100|12328_  & \new_Sorter100|12329_ ;
  assign \new_Sorter100|12429_  = \new_Sorter100|12328_  | \new_Sorter100|12329_ ;
  assign \new_Sorter100|12430_  = \new_Sorter100|12330_  & \new_Sorter100|12331_ ;
  assign \new_Sorter100|12431_  = \new_Sorter100|12330_  | \new_Sorter100|12331_ ;
  assign \new_Sorter100|12432_  = \new_Sorter100|12332_  & \new_Sorter100|12333_ ;
  assign \new_Sorter100|12433_  = \new_Sorter100|12332_  | \new_Sorter100|12333_ ;
  assign \new_Sorter100|12434_  = \new_Sorter100|12334_  & \new_Sorter100|12335_ ;
  assign \new_Sorter100|12435_  = \new_Sorter100|12334_  | \new_Sorter100|12335_ ;
  assign \new_Sorter100|12436_  = \new_Sorter100|12336_  & \new_Sorter100|12337_ ;
  assign \new_Sorter100|12437_  = \new_Sorter100|12336_  | \new_Sorter100|12337_ ;
  assign \new_Sorter100|12438_  = \new_Sorter100|12338_  & \new_Sorter100|12339_ ;
  assign \new_Sorter100|12439_  = \new_Sorter100|12338_  | \new_Sorter100|12339_ ;
  assign \new_Sorter100|12440_  = \new_Sorter100|12340_  & \new_Sorter100|12341_ ;
  assign \new_Sorter100|12441_  = \new_Sorter100|12340_  | \new_Sorter100|12341_ ;
  assign \new_Sorter100|12442_  = \new_Sorter100|12342_  & \new_Sorter100|12343_ ;
  assign \new_Sorter100|12443_  = \new_Sorter100|12342_  | \new_Sorter100|12343_ ;
  assign \new_Sorter100|12444_  = \new_Sorter100|12344_  & \new_Sorter100|12345_ ;
  assign \new_Sorter100|12445_  = \new_Sorter100|12344_  | \new_Sorter100|12345_ ;
  assign \new_Sorter100|12446_  = \new_Sorter100|12346_  & \new_Sorter100|12347_ ;
  assign \new_Sorter100|12447_  = \new_Sorter100|12346_  | \new_Sorter100|12347_ ;
  assign \new_Sorter100|12448_  = \new_Sorter100|12348_  & \new_Sorter100|12349_ ;
  assign \new_Sorter100|12449_  = \new_Sorter100|12348_  | \new_Sorter100|12349_ ;
  assign \new_Sorter100|12450_  = \new_Sorter100|12350_  & \new_Sorter100|12351_ ;
  assign \new_Sorter100|12451_  = \new_Sorter100|12350_  | \new_Sorter100|12351_ ;
  assign \new_Sorter100|12452_  = \new_Sorter100|12352_  & \new_Sorter100|12353_ ;
  assign \new_Sorter100|12453_  = \new_Sorter100|12352_  | \new_Sorter100|12353_ ;
  assign \new_Sorter100|12454_  = \new_Sorter100|12354_  & \new_Sorter100|12355_ ;
  assign \new_Sorter100|12455_  = \new_Sorter100|12354_  | \new_Sorter100|12355_ ;
  assign \new_Sorter100|12456_  = \new_Sorter100|12356_  & \new_Sorter100|12357_ ;
  assign \new_Sorter100|12457_  = \new_Sorter100|12356_  | \new_Sorter100|12357_ ;
  assign \new_Sorter100|12458_  = \new_Sorter100|12358_  & \new_Sorter100|12359_ ;
  assign \new_Sorter100|12459_  = \new_Sorter100|12358_  | \new_Sorter100|12359_ ;
  assign \new_Sorter100|12460_  = \new_Sorter100|12360_  & \new_Sorter100|12361_ ;
  assign \new_Sorter100|12461_  = \new_Sorter100|12360_  | \new_Sorter100|12361_ ;
  assign \new_Sorter100|12462_  = \new_Sorter100|12362_  & \new_Sorter100|12363_ ;
  assign \new_Sorter100|12463_  = \new_Sorter100|12362_  | \new_Sorter100|12363_ ;
  assign \new_Sorter100|12464_  = \new_Sorter100|12364_  & \new_Sorter100|12365_ ;
  assign \new_Sorter100|12465_  = \new_Sorter100|12364_  | \new_Sorter100|12365_ ;
  assign \new_Sorter100|12466_  = \new_Sorter100|12366_  & \new_Sorter100|12367_ ;
  assign \new_Sorter100|12467_  = \new_Sorter100|12366_  | \new_Sorter100|12367_ ;
  assign \new_Sorter100|12468_  = \new_Sorter100|12368_  & \new_Sorter100|12369_ ;
  assign \new_Sorter100|12469_  = \new_Sorter100|12368_  | \new_Sorter100|12369_ ;
  assign \new_Sorter100|12470_  = \new_Sorter100|12370_  & \new_Sorter100|12371_ ;
  assign \new_Sorter100|12471_  = \new_Sorter100|12370_  | \new_Sorter100|12371_ ;
  assign \new_Sorter100|12472_  = \new_Sorter100|12372_  & \new_Sorter100|12373_ ;
  assign \new_Sorter100|12473_  = \new_Sorter100|12372_  | \new_Sorter100|12373_ ;
  assign \new_Sorter100|12474_  = \new_Sorter100|12374_  & \new_Sorter100|12375_ ;
  assign \new_Sorter100|12475_  = \new_Sorter100|12374_  | \new_Sorter100|12375_ ;
  assign \new_Sorter100|12476_  = \new_Sorter100|12376_  & \new_Sorter100|12377_ ;
  assign \new_Sorter100|12477_  = \new_Sorter100|12376_  | \new_Sorter100|12377_ ;
  assign \new_Sorter100|12478_  = \new_Sorter100|12378_  & \new_Sorter100|12379_ ;
  assign \new_Sorter100|12479_  = \new_Sorter100|12378_  | \new_Sorter100|12379_ ;
  assign \new_Sorter100|12480_  = \new_Sorter100|12380_  & \new_Sorter100|12381_ ;
  assign \new_Sorter100|12481_  = \new_Sorter100|12380_  | \new_Sorter100|12381_ ;
  assign \new_Sorter100|12482_  = \new_Sorter100|12382_  & \new_Sorter100|12383_ ;
  assign \new_Sorter100|12483_  = \new_Sorter100|12382_  | \new_Sorter100|12383_ ;
  assign \new_Sorter100|12484_  = \new_Sorter100|12384_  & \new_Sorter100|12385_ ;
  assign \new_Sorter100|12485_  = \new_Sorter100|12384_  | \new_Sorter100|12385_ ;
  assign \new_Sorter100|12486_  = \new_Sorter100|12386_  & \new_Sorter100|12387_ ;
  assign \new_Sorter100|12487_  = \new_Sorter100|12386_  | \new_Sorter100|12387_ ;
  assign \new_Sorter100|12488_  = \new_Sorter100|12388_  & \new_Sorter100|12389_ ;
  assign \new_Sorter100|12489_  = \new_Sorter100|12388_  | \new_Sorter100|12389_ ;
  assign \new_Sorter100|12490_  = \new_Sorter100|12390_  & \new_Sorter100|12391_ ;
  assign \new_Sorter100|12491_  = \new_Sorter100|12390_  | \new_Sorter100|12391_ ;
  assign \new_Sorter100|12492_  = \new_Sorter100|12392_  & \new_Sorter100|12393_ ;
  assign \new_Sorter100|12493_  = \new_Sorter100|12392_  | \new_Sorter100|12393_ ;
  assign \new_Sorter100|12494_  = \new_Sorter100|12394_  & \new_Sorter100|12395_ ;
  assign \new_Sorter100|12495_  = \new_Sorter100|12394_  | \new_Sorter100|12395_ ;
  assign \new_Sorter100|12496_  = \new_Sorter100|12396_  & \new_Sorter100|12397_ ;
  assign \new_Sorter100|12497_  = \new_Sorter100|12396_  | \new_Sorter100|12397_ ;
  assign \new_Sorter100|12498_  = \new_Sorter100|12398_  & \new_Sorter100|12399_ ;
  assign \new_Sorter100|12499_  = \new_Sorter100|12398_  | \new_Sorter100|12399_ ;
  assign \new_Sorter100|12500_  = \new_Sorter100|12400_ ;
  assign \new_Sorter100|12599_  = \new_Sorter100|12499_ ;
  assign \new_Sorter100|12501_  = \new_Sorter100|12401_  & \new_Sorter100|12402_ ;
  assign \new_Sorter100|12502_  = \new_Sorter100|12401_  | \new_Sorter100|12402_ ;
  assign \new_Sorter100|12503_  = \new_Sorter100|12403_  & \new_Sorter100|12404_ ;
  assign \new_Sorter100|12504_  = \new_Sorter100|12403_  | \new_Sorter100|12404_ ;
  assign \new_Sorter100|12505_  = \new_Sorter100|12405_  & \new_Sorter100|12406_ ;
  assign \new_Sorter100|12506_  = \new_Sorter100|12405_  | \new_Sorter100|12406_ ;
  assign \new_Sorter100|12507_  = \new_Sorter100|12407_  & \new_Sorter100|12408_ ;
  assign \new_Sorter100|12508_  = \new_Sorter100|12407_  | \new_Sorter100|12408_ ;
  assign \new_Sorter100|12509_  = \new_Sorter100|12409_  & \new_Sorter100|12410_ ;
  assign \new_Sorter100|12510_  = \new_Sorter100|12409_  | \new_Sorter100|12410_ ;
  assign \new_Sorter100|12511_  = \new_Sorter100|12411_  & \new_Sorter100|12412_ ;
  assign \new_Sorter100|12512_  = \new_Sorter100|12411_  | \new_Sorter100|12412_ ;
  assign \new_Sorter100|12513_  = \new_Sorter100|12413_  & \new_Sorter100|12414_ ;
  assign \new_Sorter100|12514_  = \new_Sorter100|12413_  | \new_Sorter100|12414_ ;
  assign \new_Sorter100|12515_  = \new_Sorter100|12415_  & \new_Sorter100|12416_ ;
  assign \new_Sorter100|12516_  = \new_Sorter100|12415_  | \new_Sorter100|12416_ ;
  assign \new_Sorter100|12517_  = \new_Sorter100|12417_  & \new_Sorter100|12418_ ;
  assign \new_Sorter100|12518_  = \new_Sorter100|12417_  | \new_Sorter100|12418_ ;
  assign \new_Sorter100|12519_  = \new_Sorter100|12419_  & \new_Sorter100|12420_ ;
  assign \new_Sorter100|12520_  = \new_Sorter100|12419_  | \new_Sorter100|12420_ ;
  assign \new_Sorter100|12521_  = \new_Sorter100|12421_  & \new_Sorter100|12422_ ;
  assign \new_Sorter100|12522_  = \new_Sorter100|12421_  | \new_Sorter100|12422_ ;
  assign \new_Sorter100|12523_  = \new_Sorter100|12423_  & \new_Sorter100|12424_ ;
  assign \new_Sorter100|12524_  = \new_Sorter100|12423_  | \new_Sorter100|12424_ ;
  assign \new_Sorter100|12525_  = \new_Sorter100|12425_  & \new_Sorter100|12426_ ;
  assign \new_Sorter100|12526_  = \new_Sorter100|12425_  | \new_Sorter100|12426_ ;
  assign \new_Sorter100|12527_  = \new_Sorter100|12427_  & \new_Sorter100|12428_ ;
  assign \new_Sorter100|12528_  = \new_Sorter100|12427_  | \new_Sorter100|12428_ ;
  assign \new_Sorter100|12529_  = \new_Sorter100|12429_  & \new_Sorter100|12430_ ;
  assign \new_Sorter100|12530_  = \new_Sorter100|12429_  | \new_Sorter100|12430_ ;
  assign \new_Sorter100|12531_  = \new_Sorter100|12431_  & \new_Sorter100|12432_ ;
  assign \new_Sorter100|12532_  = \new_Sorter100|12431_  | \new_Sorter100|12432_ ;
  assign \new_Sorter100|12533_  = \new_Sorter100|12433_  & \new_Sorter100|12434_ ;
  assign \new_Sorter100|12534_  = \new_Sorter100|12433_  | \new_Sorter100|12434_ ;
  assign \new_Sorter100|12535_  = \new_Sorter100|12435_  & \new_Sorter100|12436_ ;
  assign \new_Sorter100|12536_  = \new_Sorter100|12435_  | \new_Sorter100|12436_ ;
  assign \new_Sorter100|12537_  = \new_Sorter100|12437_  & \new_Sorter100|12438_ ;
  assign \new_Sorter100|12538_  = \new_Sorter100|12437_  | \new_Sorter100|12438_ ;
  assign \new_Sorter100|12539_  = \new_Sorter100|12439_  & \new_Sorter100|12440_ ;
  assign \new_Sorter100|12540_  = \new_Sorter100|12439_  | \new_Sorter100|12440_ ;
  assign \new_Sorter100|12541_  = \new_Sorter100|12441_  & \new_Sorter100|12442_ ;
  assign \new_Sorter100|12542_  = \new_Sorter100|12441_  | \new_Sorter100|12442_ ;
  assign \new_Sorter100|12543_  = \new_Sorter100|12443_  & \new_Sorter100|12444_ ;
  assign \new_Sorter100|12544_  = \new_Sorter100|12443_  | \new_Sorter100|12444_ ;
  assign \new_Sorter100|12545_  = \new_Sorter100|12445_  & \new_Sorter100|12446_ ;
  assign \new_Sorter100|12546_  = \new_Sorter100|12445_  | \new_Sorter100|12446_ ;
  assign \new_Sorter100|12547_  = \new_Sorter100|12447_  & \new_Sorter100|12448_ ;
  assign \new_Sorter100|12548_  = \new_Sorter100|12447_  | \new_Sorter100|12448_ ;
  assign \new_Sorter100|12549_  = \new_Sorter100|12449_  & \new_Sorter100|12450_ ;
  assign \new_Sorter100|12550_  = \new_Sorter100|12449_  | \new_Sorter100|12450_ ;
  assign \new_Sorter100|12551_  = \new_Sorter100|12451_  & \new_Sorter100|12452_ ;
  assign \new_Sorter100|12552_  = \new_Sorter100|12451_  | \new_Sorter100|12452_ ;
  assign \new_Sorter100|12553_  = \new_Sorter100|12453_  & \new_Sorter100|12454_ ;
  assign \new_Sorter100|12554_  = \new_Sorter100|12453_  | \new_Sorter100|12454_ ;
  assign \new_Sorter100|12555_  = \new_Sorter100|12455_  & \new_Sorter100|12456_ ;
  assign \new_Sorter100|12556_  = \new_Sorter100|12455_  | \new_Sorter100|12456_ ;
  assign \new_Sorter100|12557_  = \new_Sorter100|12457_  & \new_Sorter100|12458_ ;
  assign \new_Sorter100|12558_  = \new_Sorter100|12457_  | \new_Sorter100|12458_ ;
  assign \new_Sorter100|12559_  = \new_Sorter100|12459_  & \new_Sorter100|12460_ ;
  assign \new_Sorter100|12560_  = \new_Sorter100|12459_  | \new_Sorter100|12460_ ;
  assign \new_Sorter100|12561_  = \new_Sorter100|12461_  & \new_Sorter100|12462_ ;
  assign \new_Sorter100|12562_  = \new_Sorter100|12461_  | \new_Sorter100|12462_ ;
  assign \new_Sorter100|12563_  = \new_Sorter100|12463_  & \new_Sorter100|12464_ ;
  assign \new_Sorter100|12564_  = \new_Sorter100|12463_  | \new_Sorter100|12464_ ;
  assign \new_Sorter100|12565_  = \new_Sorter100|12465_  & \new_Sorter100|12466_ ;
  assign \new_Sorter100|12566_  = \new_Sorter100|12465_  | \new_Sorter100|12466_ ;
  assign \new_Sorter100|12567_  = \new_Sorter100|12467_  & \new_Sorter100|12468_ ;
  assign \new_Sorter100|12568_  = \new_Sorter100|12467_  | \new_Sorter100|12468_ ;
  assign \new_Sorter100|12569_  = \new_Sorter100|12469_  & \new_Sorter100|12470_ ;
  assign \new_Sorter100|12570_  = \new_Sorter100|12469_  | \new_Sorter100|12470_ ;
  assign \new_Sorter100|12571_  = \new_Sorter100|12471_  & \new_Sorter100|12472_ ;
  assign \new_Sorter100|12572_  = \new_Sorter100|12471_  | \new_Sorter100|12472_ ;
  assign \new_Sorter100|12573_  = \new_Sorter100|12473_  & \new_Sorter100|12474_ ;
  assign \new_Sorter100|12574_  = \new_Sorter100|12473_  | \new_Sorter100|12474_ ;
  assign \new_Sorter100|12575_  = \new_Sorter100|12475_  & \new_Sorter100|12476_ ;
  assign \new_Sorter100|12576_  = \new_Sorter100|12475_  | \new_Sorter100|12476_ ;
  assign \new_Sorter100|12577_  = \new_Sorter100|12477_  & \new_Sorter100|12478_ ;
  assign \new_Sorter100|12578_  = \new_Sorter100|12477_  | \new_Sorter100|12478_ ;
  assign \new_Sorter100|12579_  = \new_Sorter100|12479_  & \new_Sorter100|12480_ ;
  assign \new_Sorter100|12580_  = \new_Sorter100|12479_  | \new_Sorter100|12480_ ;
  assign \new_Sorter100|12581_  = \new_Sorter100|12481_  & \new_Sorter100|12482_ ;
  assign \new_Sorter100|12582_  = \new_Sorter100|12481_  | \new_Sorter100|12482_ ;
  assign \new_Sorter100|12583_  = \new_Sorter100|12483_  & \new_Sorter100|12484_ ;
  assign \new_Sorter100|12584_  = \new_Sorter100|12483_  | \new_Sorter100|12484_ ;
  assign \new_Sorter100|12585_  = \new_Sorter100|12485_  & \new_Sorter100|12486_ ;
  assign \new_Sorter100|12586_  = \new_Sorter100|12485_  | \new_Sorter100|12486_ ;
  assign \new_Sorter100|12587_  = \new_Sorter100|12487_  & \new_Sorter100|12488_ ;
  assign \new_Sorter100|12588_  = \new_Sorter100|12487_  | \new_Sorter100|12488_ ;
  assign \new_Sorter100|12589_  = \new_Sorter100|12489_  & \new_Sorter100|12490_ ;
  assign \new_Sorter100|12590_  = \new_Sorter100|12489_  | \new_Sorter100|12490_ ;
  assign \new_Sorter100|12591_  = \new_Sorter100|12491_  & \new_Sorter100|12492_ ;
  assign \new_Sorter100|12592_  = \new_Sorter100|12491_  | \new_Sorter100|12492_ ;
  assign \new_Sorter100|12593_  = \new_Sorter100|12493_  & \new_Sorter100|12494_ ;
  assign \new_Sorter100|12594_  = \new_Sorter100|12493_  | \new_Sorter100|12494_ ;
  assign \new_Sorter100|12595_  = \new_Sorter100|12495_  & \new_Sorter100|12496_ ;
  assign \new_Sorter100|12596_  = \new_Sorter100|12495_  | \new_Sorter100|12496_ ;
  assign \new_Sorter100|12597_  = \new_Sorter100|12497_  & \new_Sorter100|12498_ ;
  assign \new_Sorter100|12598_  = \new_Sorter100|12497_  | \new_Sorter100|12498_ ;
  assign \new_Sorter100|12600_  = \new_Sorter100|12500_  & \new_Sorter100|12501_ ;
  assign \new_Sorter100|12601_  = \new_Sorter100|12500_  | \new_Sorter100|12501_ ;
  assign \new_Sorter100|12602_  = \new_Sorter100|12502_  & \new_Sorter100|12503_ ;
  assign \new_Sorter100|12603_  = \new_Sorter100|12502_  | \new_Sorter100|12503_ ;
  assign \new_Sorter100|12604_  = \new_Sorter100|12504_  & \new_Sorter100|12505_ ;
  assign \new_Sorter100|12605_  = \new_Sorter100|12504_  | \new_Sorter100|12505_ ;
  assign \new_Sorter100|12606_  = \new_Sorter100|12506_  & \new_Sorter100|12507_ ;
  assign \new_Sorter100|12607_  = \new_Sorter100|12506_  | \new_Sorter100|12507_ ;
  assign \new_Sorter100|12608_  = \new_Sorter100|12508_  & \new_Sorter100|12509_ ;
  assign \new_Sorter100|12609_  = \new_Sorter100|12508_  | \new_Sorter100|12509_ ;
  assign \new_Sorter100|12610_  = \new_Sorter100|12510_  & \new_Sorter100|12511_ ;
  assign \new_Sorter100|12611_  = \new_Sorter100|12510_  | \new_Sorter100|12511_ ;
  assign \new_Sorter100|12612_  = \new_Sorter100|12512_  & \new_Sorter100|12513_ ;
  assign \new_Sorter100|12613_  = \new_Sorter100|12512_  | \new_Sorter100|12513_ ;
  assign \new_Sorter100|12614_  = \new_Sorter100|12514_  & \new_Sorter100|12515_ ;
  assign \new_Sorter100|12615_  = \new_Sorter100|12514_  | \new_Sorter100|12515_ ;
  assign \new_Sorter100|12616_  = \new_Sorter100|12516_  & \new_Sorter100|12517_ ;
  assign \new_Sorter100|12617_  = \new_Sorter100|12516_  | \new_Sorter100|12517_ ;
  assign \new_Sorter100|12618_  = \new_Sorter100|12518_  & \new_Sorter100|12519_ ;
  assign \new_Sorter100|12619_  = \new_Sorter100|12518_  | \new_Sorter100|12519_ ;
  assign \new_Sorter100|12620_  = \new_Sorter100|12520_  & \new_Sorter100|12521_ ;
  assign \new_Sorter100|12621_  = \new_Sorter100|12520_  | \new_Sorter100|12521_ ;
  assign \new_Sorter100|12622_  = \new_Sorter100|12522_  & \new_Sorter100|12523_ ;
  assign \new_Sorter100|12623_  = \new_Sorter100|12522_  | \new_Sorter100|12523_ ;
  assign \new_Sorter100|12624_  = \new_Sorter100|12524_  & \new_Sorter100|12525_ ;
  assign \new_Sorter100|12625_  = \new_Sorter100|12524_  | \new_Sorter100|12525_ ;
  assign \new_Sorter100|12626_  = \new_Sorter100|12526_  & \new_Sorter100|12527_ ;
  assign \new_Sorter100|12627_  = \new_Sorter100|12526_  | \new_Sorter100|12527_ ;
  assign \new_Sorter100|12628_  = \new_Sorter100|12528_  & \new_Sorter100|12529_ ;
  assign \new_Sorter100|12629_  = \new_Sorter100|12528_  | \new_Sorter100|12529_ ;
  assign \new_Sorter100|12630_  = \new_Sorter100|12530_  & \new_Sorter100|12531_ ;
  assign \new_Sorter100|12631_  = \new_Sorter100|12530_  | \new_Sorter100|12531_ ;
  assign \new_Sorter100|12632_  = \new_Sorter100|12532_  & \new_Sorter100|12533_ ;
  assign \new_Sorter100|12633_  = \new_Sorter100|12532_  | \new_Sorter100|12533_ ;
  assign \new_Sorter100|12634_  = \new_Sorter100|12534_  & \new_Sorter100|12535_ ;
  assign \new_Sorter100|12635_  = \new_Sorter100|12534_  | \new_Sorter100|12535_ ;
  assign \new_Sorter100|12636_  = \new_Sorter100|12536_  & \new_Sorter100|12537_ ;
  assign \new_Sorter100|12637_  = \new_Sorter100|12536_  | \new_Sorter100|12537_ ;
  assign \new_Sorter100|12638_  = \new_Sorter100|12538_  & \new_Sorter100|12539_ ;
  assign \new_Sorter100|12639_  = \new_Sorter100|12538_  | \new_Sorter100|12539_ ;
  assign \new_Sorter100|12640_  = \new_Sorter100|12540_  & \new_Sorter100|12541_ ;
  assign \new_Sorter100|12641_  = \new_Sorter100|12540_  | \new_Sorter100|12541_ ;
  assign \new_Sorter100|12642_  = \new_Sorter100|12542_  & \new_Sorter100|12543_ ;
  assign \new_Sorter100|12643_  = \new_Sorter100|12542_  | \new_Sorter100|12543_ ;
  assign \new_Sorter100|12644_  = \new_Sorter100|12544_  & \new_Sorter100|12545_ ;
  assign \new_Sorter100|12645_  = \new_Sorter100|12544_  | \new_Sorter100|12545_ ;
  assign \new_Sorter100|12646_  = \new_Sorter100|12546_  & \new_Sorter100|12547_ ;
  assign \new_Sorter100|12647_  = \new_Sorter100|12546_  | \new_Sorter100|12547_ ;
  assign \new_Sorter100|12648_  = \new_Sorter100|12548_  & \new_Sorter100|12549_ ;
  assign \new_Sorter100|12649_  = \new_Sorter100|12548_  | \new_Sorter100|12549_ ;
  assign \new_Sorter100|12650_  = \new_Sorter100|12550_  & \new_Sorter100|12551_ ;
  assign \new_Sorter100|12651_  = \new_Sorter100|12550_  | \new_Sorter100|12551_ ;
  assign \new_Sorter100|12652_  = \new_Sorter100|12552_  & \new_Sorter100|12553_ ;
  assign \new_Sorter100|12653_  = \new_Sorter100|12552_  | \new_Sorter100|12553_ ;
  assign \new_Sorter100|12654_  = \new_Sorter100|12554_  & \new_Sorter100|12555_ ;
  assign \new_Sorter100|12655_  = \new_Sorter100|12554_  | \new_Sorter100|12555_ ;
  assign \new_Sorter100|12656_  = \new_Sorter100|12556_  & \new_Sorter100|12557_ ;
  assign \new_Sorter100|12657_  = \new_Sorter100|12556_  | \new_Sorter100|12557_ ;
  assign \new_Sorter100|12658_  = \new_Sorter100|12558_  & \new_Sorter100|12559_ ;
  assign \new_Sorter100|12659_  = \new_Sorter100|12558_  | \new_Sorter100|12559_ ;
  assign \new_Sorter100|12660_  = \new_Sorter100|12560_  & \new_Sorter100|12561_ ;
  assign \new_Sorter100|12661_  = \new_Sorter100|12560_  | \new_Sorter100|12561_ ;
  assign \new_Sorter100|12662_  = \new_Sorter100|12562_  & \new_Sorter100|12563_ ;
  assign \new_Sorter100|12663_  = \new_Sorter100|12562_  | \new_Sorter100|12563_ ;
  assign \new_Sorter100|12664_  = \new_Sorter100|12564_  & \new_Sorter100|12565_ ;
  assign \new_Sorter100|12665_  = \new_Sorter100|12564_  | \new_Sorter100|12565_ ;
  assign \new_Sorter100|12666_  = \new_Sorter100|12566_  & \new_Sorter100|12567_ ;
  assign \new_Sorter100|12667_  = \new_Sorter100|12566_  | \new_Sorter100|12567_ ;
  assign \new_Sorter100|12668_  = \new_Sorter100|12568_  & \new_Sorter100|12569_ ;
  assign \new_Sorter100|12669_  = \new_Sorter100|12568_  | \new_Sorter100|12569_ ;
  assign \new_Sorter100|12670_  = \new_Sorter100|12570_  & \new_Sorter100|12571_ ;
  assign \new_Sorter100|12671_  = \new_Sorter100|12570_  | \new_Sorter100|12571_ ;
  assign \new_Sorter100|12672_  = \new_Sorter100|12572_  & \new_Sorter100|12573_ ;
  assign \new_Sorter100|12673_  = \new_Sorter100|12572_  | \new_Sorter100|12573_ ;
  assign \new_Sorter100|12674_  = \new_Sorter100|12574_  & \new_Sorter100|12575_ ;
  assign \new_Sorter100|12675_  = \new_Sorter100|12574_  | \new_Sorter100|12575_ ;
  assign \new_Sorter100|12676_  = \new_Sorter100|12576_  & \new_Sorter100|12577_ ;
  assign \new_Sorter100|12677_  = \new_Sorter100|12576_  | \new_Sorter100|12577_ ;
  assign \new_Sorter100|12678_  = \new_Sorter100|12578_  & \new_Sorter100|12579_ ;
  assign \new_Sorter100|12679_  = \new_Sorter100|12578_  | \new_Sorter100|12579_ ;
  assign \new_Sorter100|12680_  = \new_Sorter100|12580_  & \new_Sorter100|12581_ ;
  assign \new_Sorter100|12681_  = \new_Sorter100|12580_  | \new_Sorter100|12581_ ;
  assign \new_Sorter100|12682_  = \new_Sorter100|12582_  & \new_Sorter100|12583_ ;
  assign \new_Sorter100|12683_  = \new_Sorter100|12582_  | \new_Sorter100|12583_ ;
  assign \new_Sorter100|12684_  = \new_Sorter100|12584_  & \new_Sorter100|12585_ ;
  assign \new_Sorter100|12685_  = \new_Sorter100|12584_  | \new_Sorter100|12585_ ;
  assign \new_Sorter100|12686_  = \new_Sorter100|12586_  & \new_Sorter100|12587_ ;
  assign \new_Sorter100|12687_  = \new_Sorter100|12586_  | \new_Sorter100|12587_ ;
  assign \new_Sorter100|12688_  = \new_Sorter100|12588_  & \new_Sorter100|12589_ ;
  assign \new_Sorter100|12689_  = \new_Sorter100|12588_  | \new_Sorter100|12589_ ;
  assign \new_Sorter100|12690_  = \new_Sorter100|12590_  & \new_Sorter100|12591_ ;
  assign \new_Sorter100|12691_  = \new_Sorter100|12590_  | \new_Sorter100|12591_ ;
  assign \new_Sorter100|12692_  = \new_Sorter100|12592_  & \new_Sorter100|12593_ ;
  assign \new_Sorter100|12693_  = \new_Sorter100|12592_  | \new_Sorter100|12593_ ;
  assign \new_Sorter100|12694_  = \new_Sorter100|12594_  & \new_Sorter100|12595_ ;
  assign \new_Sorter100|12695_  = \new_Sorter100|12594_  | \new_Sorter100|12595_ ;
  assign \new_Sorter100|12696_  = \new_Sorter100|12596_  & \new_Sorter100|12597_ ;
  assign \new_Sorter100|12697_  = \new_Sorter100|12596_  | \new_Sorter100|12597_ ;
  assign \new_Sorter100|12698_  = \new_Sorter100|12598_  & \new_Sorter100|12599_ ;
  assign \new_Sorter100|12699_  = \new_Sorter100|12598_  | \new_Sorter100|12599_ ;
  assign \new_Sorter100|12700_  = \new_Sorter100|12600_ ;
  assign \new_Sorter100|12799_  = \new_Sorter100|12699_ ;
  assign \new_Sorter100|12701_  = \new_Sorter100|12601_  & \new_Sorter100|12602_ ;
  assign \new_Sorter100|12702_  = \new_Sorter100|12601_  | \new_Sorter100|12602_ ;
  assign \new_Sorter100|12703_  = \new_Sorter100|12603_  & \new_Sorter100|12604_ ;
  assign \new_Sorter100|12704_  = \new_Sorter100|12603_  | \new_Sorter100|12604_ ;
  assign \new_Sorter100|12705_  = \new_Sorter100|12605_  & \new_Sorter100|12606_ ;
  assign \new_Sorter100|12706_  = \new_Sorter100|12605_  | \new_Sorter100|12606_ ;
  assign \new_Sorter100|12707_  = \new_Sorter100|12607_  & \new_Sorter100|12608_ ;
  assign \new_Sorter100|12708_  = \new_Sorter100|12607_  | \new_Sorter100|12608_ ;
  assign \new_Sorter100|12709_  = \new_Sorter100|12609_  & \new_Sorter100|12610_ ;
  assign \new_Sorter100|12710_  = \new_Sorter100|12609_  | \new_Sorter100|12610_ ;
  assign \new_Sorter100|12711_  = \new_Sorter100|12611_  & \new_Sorter100|12612_ ;
  assign \new_Sorter100|12712_  = \new_Sorter100|12611_  | \new_Sorter100|12612_ ;
  assign \new_Sorter100|12713_  = \new_Sorter100|12613_  & \new_Sorter100|12614_ ;
  assign \new_Sorter100|12714_  = \new_Sorter100|12613_  | \new_Sorter100|12614_ ;
  assign \new_Sorter100|12715_  = \new_Sorter100|12615_  & \new_Sorter100|12616_ ;
  assign \new_Sorter100|12716_  = \new_Sorter100|12615_  | \new_Sorter100|12616_ ;
  assign \new_Sorter100|12717_  = \new_Sorter100|12617_  & \new_Sorter100|12618_ ;
  assign \new_Sorter100|12718_  = \new_Sorter100|12617_  | \new_Sorter100|12618_ ;
  assign \new_Sorter100|12719_  = \new_Sorter100|12619_  & \new_Sorter100|12620_ ;
  assign \new_Sorter100|12720_  = \new_Sorter100|12619_  | \new_Sorter100|12620_ ;
  assign \new_Sorter100|12721_  = \new_Sorter100|12621_  & \new_Sorter100|12622_ ;
  assign \new_Sorter100|12722_  = \new_Sorter100|12621_  | \new_Sorter100|12622_ ;
  assign \new_Sorter100|12723_  = \new_Sorter100|12623_  & \new_Sorter100|12624_ ;
  assign \new_Sorter100|12724_  = \new_Sorter100|12623_  | \new_Sorter100|12624_ ;
  assign \new_Sorter100|12725_  = \new_Sorter100|12625_  & \new_Sorter100|12626_ ;
  assign \new_Sorter100|12726_  = \new_Sorter100|12625_  | \new_Sorter100|12626_ ;
  assign \new_Sorter100|12727_  = \new_Sorter100|12627_  & \new_Sorter100|12628_ ;
  assign \new_Sorter100|12728_  = \new_Sorter100|12627_  | \new_Sorter100|12628_ ;
  assign \new_Sorter100|12729_  = \new_Sorter100|12629_  & \new_Sorter100|12630_ ;
  assign \new_Sorter100|12730_  = \new_Sorter100|12629_  | \new_Sorter100|12630_ ;
  assign \new_Sorter100|12731_  = \new_Sorter100|12631_  & \new_Sorter100|12632_ ;
  assign \new_Sorter100|12732_  = \new_Sorter100|12631_  | \new_Sorter100|12632_ ;
  assign \new_Sorter100|12733_  = \new_Sorter100|12633_  & \new_Sorter100|12634_ ;
  assign \new_Sorter100|12734_  = \new_Sorter100|12633_  | \new_Sorter100|12634_ ;
  assign \new_Sorter100|12735_  = \new_Sorter100|12635_  & \new_Sorter100|12636_ ;
  assign \new_Sorter100|12736_  = \new_Sorter100|12635_  | \new_Sorter100|12636_ ;
  assign \new_Sorter100|12737_  = \new_Sorter100|12637_  & \new_Sorter100|12638_ ;
  assign \new_Sorter100|12738_  = \new_Sorter100|12637_  | \new_Sorter100|12638_ ;
  assign \new_Sorter100|12739_  = \new_Sorter100|12639_  & \new_Sorter100|12640_ ;
  assign \new_Sorter100|12740_  = \new_Sorter100|12639_  | \new_Sorter100|12640_ ;
  assign \new_Sorter100|12741_  = \new_Sorter100|12641_  & \new_Sorter100|12642_ ;
  assign \new_Sorter100|12742_  = \new_Sorter100|12641_  | \new_Sorter100|12642_ ;
  assign \new_Sorter100|12743_  = \new_Sorter100|12643_  & \new_Sorter100|12644_ ;
  assign \new_Sorter100|12744_  = \new_Sorter100|12643_  | \new_Sorter100|12644_ ;
  assign \new_Sorter100|12745_  = \new_Sorter100|12645_  & \new_Sorter100|12646_ ;
  assign \new_Sorter100|12746_  = \new_Sorter100|12645_  | \new_Sorter100|12646_ ;
  assign \new_Sorter100|12747_  = \new_Sorter100|12647_  & \new_Sorter100|12648_ ;
  assign \new_Sorter100|12748_  = \new_Sorter100|12647_  | \new_Sorter100|12648_ ;
  assign \new_Sorter100|12749_  = \new_Sorter100|12649_  & \new_Sorter100|12650_ ;
  assign \new_Sorter100|12750_  = \new_Sorter100|12649_  | \new_Sorter100|12650_ ;
  assign \new_Sorter100|12751_  = \new_Sorter100|12651_  & \new_Sorter100|12652_ ;
  assign \new_Sorter100|12752_  = \new_Sorter100|12651_  | \new_Sorter100|12652_ ;
  assign \new_Sorter100|12753_  = \new_Sorter100|12653_  & \new_Sorter100|12654_ ;
  assign \new_Sorter100|12754_  = \new_Sorter100|12653_  | \new_Sorter100|12654_ ;
  assign \new_Sorter100|12755_  = \new_Sorter100|12655_  & \new_Sorter100|12656_ ;
  assign \new_Sorter100|12756_  = \new_Sorter100|12655_  | \new_Sorter100|12656_ ;
  assign \new_Sorter100|12757_  = \new_Sorter100|12657_  & \new_Sorter100|12658_ ;
  assign \new_Sorter100|12758_  = \new_Sorter100|12657_  | \new_Sorter100|12658_ ;
  assign \new_Sorter100|12759_  = \new_Sorter100|12659_  & \new_Sorter100|12660_ ;
  assign \new_Sorter100|12760_  = \new_Sorter100|12659_  | \new_Sorter100|12660_ ;
  assign \new_Sorter100|12761_  = \new_Sorter100|12661_  & \new_Sorter100|12662_ ;
  assign \new_Sorter100|12762_  = \new_Sorter100|12661_  | \new_Sorter100|12662_ ;
  assign \new_Sorter100|12763_  = \new_Sorter100|12663_  & \new_Sorter100|12664_ ;
  assign \new_Sorter100|12764_  = \new_Sorter100|12663_  | \new_Sorter100|12664_ ;
  assign \new_Sorter100|12765_  = \new_Sorter100|12665_  & \new_Sorter100|12666_ ;
  assign \new_Sorter100|12766_  = \new_Sorter100|12665_  | \new_Sorter100|12666_ ;
  assign \new_Sorter100|12767_  = \new_Sorter100|12667_  & \new_Sorter100|12668_ ;
  assign \new_Sorter100|12768_  = \new_Sorter100|12667_  | \new_Sorter100|12668_ ;
  assign \new_Sorter100|12769_  = \new_Sorter100|12669_  & \new_Sorter100|12670_ ;
  assign \new_Sorter100|12770_  = \new_Sorter100|12669_  | \new_Sorter100|12670_ ;
  assign \new_Sorter100|12771_  = \new_Sorter100|12671_  & \new_Sorter100|12672_ ;
  assign \new_Sorter100|12772_  = \new_Sorter100|12671_  | \new_Sorter100|12672_ ;
  assign \new_Sorter100|12773_  = \new_Sorter100|12673_  & \new_Sorter100|12674_ ;
  assign \new_Sorter100|12774_  = \new_Sorter100|12673_  | \new_Sorter100|12674_ ;
  assign \new_Sorter100|12775_  = \new_Sorter100|12675_  & \new_Sorter100|12676_ ;
  assign \new_Sorter100|12776_  = \new_Sorter100|12675_  | \new_Sorter100|12676_ ;
  assign \new_Sorter100|12777_  = \new_Sorter100|12677_  & \new_Sorter100|12678_ ;
  assign \new_Sorter100|12778_  = \new_Sorter100|12677_  | \new_Sorter100|12678_ ;
  assign \new_Sorter100|12779_  = \new_Sorter100|12679_  & \new_Sorter100|12680_ ;
  assign \new_Sorter100|12780_  = \new_Sorter100|12679_  | \new_Sorter100|12680_ ;
  assign \new_Sorter100|12781_  = \new_Sorter100|12681_  & \new_Sorter100|12682_ ;
  assign \new_Sorter100|12782_  = \new_Sorter100|12681_  | \new_Sorter100|12682_ ;
  assign \new_Sorter100|12783_  = \new_Sorter100|12683_  & \new_Sorter100|12684_ ;
  assign \new_Sorter100|12784_  = \new_Sorter100|12683_  | \new_Sorter100|12684_ ;
  assign \new_Sorter100|12785_  = \new_Sorter100|12685_  & \new_Sorter100|12686_ ;
  assign \new_Sorter100|12786_  = \new_Sorter100|12685_  | \new_Sorter100|12686_ ;
  assign \new_Sorter100|12787_  = \new_Sorter100|12687_  & \new_Sorter100|12688_ ;
  assign \new_Sorter100|12788_  = \new_Sorter100|12687_  | \new_Sorter100|12688_ ;
  assign \new_Sorter100|12789_  = \new_Sorter100|12689_  & \new_Sorter100|12690_ ;
  assign \new_Sorter100|12790_  = \new_Sorter100|12689_  | \new_Sorter100|12690_ ;
  assign \new_Sorter100|12791_  = \new_Sorter100|12691_  & \new_Sorter100|12692_ ;
  assign \new_Sorter100|12792_  = \new_Sorter100|12691_  | \new_Sorter100|12692_ ;
  assign \new_Sorter100|12793_  = \new_Sorter100|12693_  & \new_Sorter100|12694_ ;
  assign \new_Sorter100|12794_  = \new_Sorter100|12693_  | \new_Sorter100|12694_ ;
  assign \new_Sorter100|12795_  = \new_Sorter100|12695_  & \new_Sorter100|12696_ ;
  assign \new_Sorter100|12796_  = \new_Sorter100|12695_  | \new_Sorter100|12696_ ;
  assign \new_Sorter100|12797_  = \new_Sorter100|12697_  & \new_Sorter100|12698_ ;
  assign \new_Sorter100|12798_  = \new_Sorter100|12697_  | \new_Sorter100|12698_ ;
  assign \new_Sorter100|12800_  = \new_Sorter100|12700_  & \new_Sorter100|12701_ ;
  assign \new_Sorter100|12801_  = \new_Sorter100|12700_  | \new_Sorter100|12701_ ;
  assign \new_Sorter100|12802_  = \new_Sorter100|12702_  & \new_Sorter100|12703_ ;
  assign \new_Sorter100|12803_  = \new_Sorter100|12702_  | \new_Sorter100|12703_ ;
  assign \new_Sorter100|12804_  = \new_Sorter100|12704_  & \new_Sorter100|12705_ ;
  assign \new_Sorter100|12805_  = \new_Sorter100|12704_  | \new_Sorter100|12705_ ;
  assign \new_Sorter100|12806_  = \new_Sorter100|12706_  & \new_Sorter100|12707_ ;
  assign \new_Sorter100|12807_  = \new_Sorter100|12706_  | \new_Sorter100|12707_ ;
  assign \new_Sorter100|12808_  = \new_Sorter100|12708_  & \new_Sorter100|12709_ ;
  assign \new_Sorter100|12809_  = \new_Sorter100|12708_  | \new_Sorter100|12709_ ;
  assign \new_Sorter100|12810_  = \new_Sorter100|12710_  & \new_Sorter100|12711_ ;
  assign \new_Sorter100|12811_  = \new_Sorter100|12710_  | \new_Sorter100|12711_ ;
  assign \new_Sorter100|12812_  = \new_Sorter100|12712_  & \new_Sorter100|12713_ ;
  assign \new_Sorter100|12813_  = \new_Sorter100|12712_  | \new_Sorter100|12713_ ;
  assign \new_Sorter100|12814_  = \new_Sorter100|12714_  & \new_Sorter100|12715_ ;
  assign \new_Sorter100|12815_  = \new_Sorter100|12714_  | \new_Sorter100|12715_ ;
  assign \new_Sorter100|12816_  = \new_Sorter100|12716_  & \new_Sorter100|12717_ ;
  assign \new_Sorter100|12817_  = \new_Sorter100|12716_  | \new_Sorter100|12717_ ;
  assign \new_Sorter100|12818_  = \new_Sorter100|12718_  & \new_Sorter100|12719_ ;
  assign \new_Sorter100|12819_  = \new_Sorter100|12718_  | \new_Sorter100|12719_ ;
  assign \new_Sorter100|12820_  = \new_Sorter100|12720_  & \new_Sorter100|12721_ ;
  assign \new_Sorter100|12821_  = \new_Sorter100|12720_  | \new_Sorter100|12721_ ;
  assign \new_Sorter100|12822_  = \new_Sorter100|12722_  & \new_Sorter100|12723_ ;
  assign \new_Sorter100|12823_  = \new_Sorter100|12722_  | \new_Sorter100|12723_ ;
  assign \new_Sorter100|12824_  = \new_Sorter100|12724_  & \new_Sorter100|12725_ ;
  assign \new_Sorter100|12825_  = \new_Sorter100|12724_  | \new_Sorter100|12725_ ;
  assign \new_Sorter100|12826_  = \new_Sorter100|12726_  & \new_Sorter100|12727_ ;
  assign \new_Sorter100|12827_  = \new_Sorter100|12726_  | \new_Sorter100|12727_ ;
  assign \new_Sorter100|12828_  = \new_Sorter100|12728_  & \new_Sorter100|12729_ ;
  assign \new_Sorter100|12829_  = \new_Sorter100|12728_  | \new_Sorter100|12729_ ;
  assign \new_Sorter100|12830_  = \new_Sorter100|12730_  & \new_Sorter100|12731_ ;
  assign \new_Sorter100|12831_  = \new_Sorter100|12730_  | \new_Sorter100|12731_ ;
  assign \new_Sorter100|12832_  = \new_Sorter100|12732_  & \new_Sorter100|12733_ ;
  assign \new_Sorter100|12833_  = \new_Sorter100|12732_  | \new_Sorter100|12733_ ;
  assign \new_Sorter100|12834_  = \new_Sorter100|12734_  & \new_Sorter100|12735_ ;
  assign \new_Sorter100|12835_  = \new_Sorter100|12734_  | \new_Sorter100|12735_ ;
  assign \new_Sorter100|12836_  = \new_Sorter100|12736_  & \new_Sorter100|12737_ ;
  assign \new_Sorter100|12837_  = \new_Sorter100|12736_  | \new_Sorter100|12737_ ;
  assign \new_Sorter100|12838_  = \new_Sorter100|12738_  & \new_Sorter100|12739_ ;
  assign \new_Sorter100|12839_  = \new_Sorter100|12738_  | \new_Sorter100|12739_ ;
  assign \new_Sorter100|12840_  = \new_Sorter100|12740_  & \new_Sorter100|12741_ ;
  assign \new_Sorter100|12841_  = \new_Sorter100|12740_  | \new_Sorter100|12741_ ;
  assign \new_Sorter100|12842_  = \new_Sorter100|12742_  & \new_Sorter100|12743_ ;
  assign \new_Sorter100|12843_  = \new_Sorter100|12742_  | \new_Sorter100|12743_ ;
  assign \new_Sorter100|12844_  = \new_Sorter100|12744_  & \new_Sorter100|12745_ ;
  assign \new_Sorter100|12845_  = \new_Sorter100|12744_  | \new_Sorter100|12745_ ;
  assign \new_Sorter100|12846_  = \new_Sorter100|12746_  & \new_Sorter100|12747_ ;
  assign \new_Sorter100|12847_  = \new_Sorter100|12746_  | \new_Sorter100|12747_ ;
  assign \new_Sorter100|12848_  = \new_Sorter100|12748_  & \new_Sorter100|12749_ ;
  assign \new_Sorter100|12849_  = \new_Sorter100|12748_  | \new_Sorter100|12749_ ;
  assign \new_Sorter100|12850_  = \new_Sorter100|12750_  & \new_Sorter100|12751_ ;
  assign \new_Sorter100|12851_  = \new_Sorter100|12750_  | \new_Sorter100|12751_ ;
  assign \new_Sorter100|12852_  = \new_Sorter100|12752_  & \new_Sorter100|12753_ ;
  assign \new_Sorter100|12853_  = \new_Sorter100|12752_  | \new_Sorter100|12753_ ;
  assign \new_Sorter100|12854_  = \new_Sorter100|12754_  & \new_Sorter100|12755_ ;
  assign \new_Sorter100|12855_  = \new_Sorter100|12754_  | \new_Sorter100|12755_ ;
  assign \new_Sorter100|12856_  = \new_Sorter100|12756_  & \new_Sorter100|12757_ ;
  assign \new_Sorter100|12857_  = \new_Sorter100|12756_  | \new_Sorter100|12757_ ;
  assign \new_Sorter100|12858_  = \new_Sorter100|12758_  & \new_Sorter100|12759_ ;
  assign \new_Sorter100|12859_  = \new_Sorter100|12758_  | \new_Sorter100|12759_ ;
  assign \new_Sorter100|12860_  = \new_Sorter100|12760_  & \new_Sorter100|12761_ ;
  assign \new_Sorter100|12861_  = \new_Sorter100|12760_  | \new_Sorter100|12761_ ;
  assign \new_Sorter100|12862_  = \new_Sorter100|12762_  & \new_Sorter100|12763_ ;
  assign \new_Sorter100|12863_  = \new_Sorter100|12762_  | \new_Sorter100|12763_ ;
  assign \new_Sorter100|12864_  = \new_Sorter100|12764_  & \new_Sorter100|12765_ ;
  assign \new_Sorter100|12865_  = \new_Sorter100|12764_  | \new_Sorter100|12765_ ;
  assign \new_Sorter100|12866_  = \new_Sorter100|12766_  & \new_Sorter100|12767_ ;
  assign \new_Sorter100|12867_  = \new_Sorter100|12766_  | \new_Sorter100|12767_ ;
  assign \new_Sorter100|12868_  = \new_Sorter100|12768_  & \new_Sorter100|12769_ ;
  assign \new_Sorter100|12869_  = \new_Sorter100|12768_  | \new_Sorter100|12769_ ;
  assign \new_Sorter100|12870_  = \new_Sorter100|12770_  & \new_Sorter100|12771_ ;
  assign \new_Sorter100|12871_  = \new_Sorter100|12770_  | \new_Sorter100|12771_ ;
  assign \new_Sorter100|12872_  = \new_Sorter100|12772_  & \new_Sorter100|12773_ ;
  assign \new_Sorter100|12873_  = \new_Sorter100|12772_  | \new_Sorter100|12773_ ;
  assign \new_Sorter100|12874_  = \new_Sorter100|12774_  & \new_Sorter100|12775_ ;
  assign \new_Sorter100|12875_  = \new_Sorter100|12774_  | \new_Sorter100|12775_ ;
  assign \new_Sorter100|12876_  = \new_Sorter100|12776_  & \new_Sorter100|12777_ ;
  assign \new_Sorter100|12877_  = \new_Sorter100|12776_  | \new_Sorter100|12777_ ;
  assign \new_Sorter100|12878_  = \new_Sorter100|12778_  & \new_Sorter100|12779_ ;
  assign \new_Sorter100|12879_  = \new_Sorter100|12778_  | \new_Sorter100|12779_ ;
  assign \new_Sorter100|12880_  = \new_Sorter100|12780_  & \new_Sorter100|12781_ ;
  assign \new_Sorter100|12881_  = \new_Sorter100|12780_  | \new_Sorter100|12781_ ;
  assign \new_Sorter100|12882_  = \new_Sorter100|12782_  & \new_Sorter100|12783_ ;
  assign \new_Sorter100|12883_  = \new_Sorter100|12782_  | \new_Sorter100|12783_ ;
  assign \new_Sorter100|12884_  = \new_Sorter100|12784_  & \new_Sorter100|12785_ ;
  assign \new_Sorter100|12885_  = \new_Sorter100|12784_  | \new_Sorter100|12785_ ;
  assign \new_Sorter100|12886_  = \new_Sorter100|12786_  & \new_Sorter100|12787_ ;
  assign \new_Sorter100|12887_  = \new_Sorter100|12786_  | \new_Sorter100|12787_ ;
  assign \new_Sorter100|12888_  = \new_Sorter100|12788_  & \new_Sorter100|12789_ ;
  assign \new_Sorter100|12889_  = \new_Sorter100|12788_  | \new_Sorter100|12789_ ;
  assign \new_Sorter100|12890_  = \new_Sorter100|12790_  & \new_Sorter100|12791_ ;
  assign \new_Sorter100|12891_  = \new_Sorter100|12790_  | \new_Sorter100|12791_ ;
  assign \new_Sorter100|12892_  = \new_Sorter100|12792_  & \new_Sorter100|12793_ ;
  assign \new_Sorter100|12893_  = \new_Sorter100|12792_  | \new_Sorter100|12793_ ;
  assign \new_Sorter100|12894_  = \new_Sorter100|12794_  & \new_Sorter100|12795_ ;
  assign \new_Sorter100|12895_  = \new_Sorter100|12794_  | \new_Sorter100|12795_ ;
  assign \new_Sorter100|12896_  = \new_Sorter100|12796_  & \new_Sorter100|12797_ ;
  assign \new_Sorter100|12897_  = \new_Sorter100|12796_  | \new_Sorter100|12797_ ;
  assign \new_Sorter100|12898_  = \new_Sorter100|12798_  & \new_Sorter100|12799_ ;
  assign \new_Sorter100|12899_  = \new_Sorter100|12798_  | \new_Sorter100|12799_ ;
  assign \new_Sorter100|12900_  = \new_Sorter100|12800_ ;
  assign \new_Sorter100|12999_  = \new_Sorter100|12899_ ;
  assign \new_Sorter100|12901_  = \new_Sorter100|12801_  & \new_Sorter100|12802_ ;
  assign \new_Sorter100|12902_  = \new_Sorter100|12801_  | \new_Sorter100|12802_ ;
  assign \new_Sorter100|12903_  = \new_Sorter100|12803_  & \new_Sorter100|12804_ ;
  assign \new_Sorter100|12904_  = \new_Sorter100|12803_  | \new_Sorter100|12804_ ;
  assign \new_Sorter100|12905_  = \new_Sorter100|12805_  & \new_Sorter100|12806_ ;
  assign \new_Sorter100|12906_  = \new_Sorter100|12805_  | \new_Sorter100|12806_ ;
  assign \new_Sorter100|12907_  = \new_Sorter100|12807_  & \new_Sorter100|12808_ ;
  assign \new_Sorter100|12908_  = \new_Sorter100|12807_  | \new_Sorter100|12808_ ;
  assign \new_Sorter100|12909_  = \new_Sorter100|12809_  & \new_Sorter100|12810_ ;
  assign \new_Sorter100|12910_  = \new_Sorter100|12809_  | \new_Sorter100|12810_ ;
  assign \new_Sorter100|12911_  = \new_Sorter100|12811_  & \new_Sorter100|12812_ ;
  assign \new_Sorter100|12912_  = \new_Sorter100|12811_  | \new_Sorter100|12812_ ;
  assign \new_Sorter100|12913_  = \new_Sorter100|12813_  & \new_Sorter100|12814_ ;
  assign \new_Sorter100|12914_  = \new_Sorter100|12813_  | \new_Sorter100|12814_ ;
  assign \new_Sorter100|12915_  = \new_Sorter100|12815_  & \new_Sorter100|12816_ ;
  assign \new_Sorter100|12916_  = \new_Sorter100|12815_  | \new_Sorter100|12816_ ;
  assign \new_Sorter100|12917_  = \new_Sorter100|12817_  & \new_Sorter100|12818_ ;
  assign \new_Sorter100|12918_  = \new_Sorter100|12817_  | \new_Sorter100|12818_ ;
  assign \new_Sorter100|12919_  = \new_Sorter100|12819_  & \new_Sorter100|12820_ ;
  assign \new_Sorter100|12920_  = \new_Sorter100|12819_  | \new_Sorter100|12820_ ;
  assign \new_Sorter100|12921_  = \new_Sorter100|12821_  & \new_Sorter100|12822_ ;
  assign \new_Sorter100|12922_  = \new_Sorter100|12821_  | \new_Sorter100|12822_ ;
  assign \new_Sorter100|12923_  = \new_Sorter100|12823_  & \new_Sorter100|12824_ ;
  assign \new_Sorter100|12924_  = \new_Sorter100|12823_  | \new_Sorter100|12824_ ;
  assign \new_Sorter100|12925_  = \new_Sorter100|12825_  & \new_Sorter100|12826_ ;
  assign \new_Sorter100|12926_  = \new_Sorter100|12825_  | \new_Sorter100|12826_ ;
  assign \new_Sorter100|12927_  = \new_Sorter100|12827_  & \new_Sorter100|12828_ ;
  assign \new_Sorter100|12928_  = \new_Sorter100|12827_  | \new_Sorter100|12828_ ;
  assign \new_Sorter100|12929_  = \new_Sorter100|12829_  & \new_Sorter100|12830_ ;
  assign \new_Sorter100|12930_  = \new_Sorter100|12829_  | \new_Sorter100|12830_ ;
  assign \new_Sorter100|12931_  = \new_Sorter100|12831_  & \new_Sorter100|12832_ ;
  assign \new_Sorter100|12932_  = \new_Sorter100|12831_  | \new_Sorter100|12832_ ;
  assign \new_Sorter100|12933_  = \new_Sorter100|12833_  & \new_Sorter100|12834_ ;
  assign \new_Sorter100|12934_  = \new_Sorter100|12833_  | \new_Sorter100|12834_ ;
  assign \new_Sorter100|12935_  = \new_Sorter100|12835_  & \new_Sorter100|12836_ ;
  assign \new_Sorter100|12936_  = \new_Sorter100|12835_  | \new_Sorter100|12836_ ;
  assign \new_Sorter100|12937_  = \new_Sorter100|12837_  & \new_Sorter100|12838_ ;
  assign \new_Sorter100|12938_  = \new_Sorter100|12837_  | \new_Sorter100|12838_ ;
  assign \new_Sorter100|12939_  = \new_Sorter100|12839_  & \new_Sorter100|12840_ ;
  assign \new_Sorter100|12940_  = \new_Sorter100|12839_  | \new_Sorter100|12840_ ;
  assign \new_Sorter100|12941_  = \new_Sorter100|12841_  & \new_Sorter100|12842_ ;
  assign \new_Sorter100|12942_  = \new_Sorter100|12841_  | \new_Sorter100|12842_ ;
  assign \new_Sorter100|12943_  = \new_Sorter100|12843_  & \new_Sorter100|12844_ ;
  assign \new_Sorter100|12944_  = \new_Sorter100|12843_  | \new_Sorter100|12844_ ;
  assign \new_Sorter100|12945_  = \new_Sorter100|12845_  & \new_Sorter100|12846_ ;
  assign \new_Sorter100|12946_  = \new_Sorter100|12845_  | \new_Sorter100|12846_ ;
  assign \new_Sorter100|12947_  = \new_Sorter100|12847_  & \new_Sorter100|12848_ ;
  assign \new_Sorter100|12948_  = \new_Sorter100|12847_  | \new_Sorter100|12848_ ;
  assign \new_Sorter100|12949_  = \new_Sorter100|12849_  & \new_Sorter100|12850_ ;
  assign \new_Sorter100|12950_  = \new_Sorter100|12849_  | \new_Sorter100|12850_ ;
  assign \new_Sorter100|12951_  = \new_Sorter100|12851_  & \new_Sorter100|12852_ ;
  assign \new_Sorter100|12952_  = \new_Sorter100|12851_  | \new_Sorter100|12852_ ;
  assign \new_Sorter100|12953_  = \new_Sorter100|12853_  & \new_Sorter100|12854_ ;
  assign \new_Sorter100|12954_  = \new_Sorter100|12853_  | \new_Sorter100|12854_ ;
  assign \new_Sorter100|12955_  = \new_Sorter100|12855_  & \new_Sorter100|12856_ ;
  assign \new_Sorter100|12956_  = \new_Sorter100|12855_  | \new_Sorter100|12856_ ;
  assign \new_Sorter100|12957_  = \new_Sorter100|12857_  & \new_Sorter100|12858_ ;
  assign \new_Sorter100|12958_  = \new_Sorter100|12857_  | \new_Sorter100|12858_ ;
  assign \new_Sorter100|12959_  = \new_Sorter100|12859_  & \new_Sorter100|12860_ ;
  assign \new_Sorter100|12960_  = \new_Sorter100|12859_  | \new_Sorter100|12860_ ;
  assign \new_Sorter100|12961_  = \new_Sorter100|12861_  & \new_Sorter100|12862_ ;
  assign \new_Sorter100|12962_  = \new_Sorter100|12861_  | \new_Sorter100|12862_ ;
  assign \new_Sorter100|12963_  = \new_Sorter100|12863_  & \new_Sorter100|12864_ ;
  assign \new_Sorter100|12964_  = \new_Sorter100|12863_  | \new_Sorter100|12864_ ;
  assign \new_Sorter100|12965_  = \new_Sorter100|12865_  & \new_Sorter100|12866_ ;
  assign \new_Sorter100|12966_  = \new_Sorter100|12865_  | \new_Sorter100|12866_ ;
  assign \new_Sorter100|12967_  = \new_Sorter100|12867_  & \new_Sorter100|12868_ ;
  assign \new_Sorter100|12968_  = \new_Sorter100|12867_  | \new_Sorter100|12868_ ;
  assign \new_Sorter100|12969_  = \new_Sorter100|12869_  & \new_Sorter100|12870_ ;
  assign \new_Sorter100|12970_  = \new_Sorter100|12869_  | \new_Sorter100|12870_ ;
  assign \new_Sorter100|12971_  = \new_Sorter100|12871_  & \new_Sorter100|12872_ ;
  assign \new_Sorter100|12972_  = \new_Sorter100|12871_  | \new_Sorter100|12872_ ;
  assign \new_Sorter100|12973_  = \new_Sorter100|12873_  & \new_Sorter100|12874_ ;
  assign \new_Sorter100|12974_  = \new_Sorter100|12873_  | \new_Sorter100|12874_ ;
  assign \new_Sorter100|12975_  = \new_Sorter100|12875_  & \new_Sorter100|12876_ ;
  assign \new_Sorter100|12976_  = \new_Sorter100|12875_  | \new_Sorter100|12876_ ;
  assign \new_Sorter100|12977_  = \new_Sorter100|12877_  & \new_Sorter100|12878_ ;
  assign \new_Sorter100|12978_  = \new_Sorter100|12877_  | \new_Sorter100|12878_ ;
  assign \new_Sorter100|12979_  = \new_Sorter100|12879_  & \new_Sorter100|12880_ ;
  assign \new_Sorter100|12980_  = \new_Sorter100|12879_  | \new_Sorter100|12880_ ;
  assign \new_Sorter100|12981_  = \new_Sorter100|12881_  & \new_Sorter100|12882_ ;
  assign \new_Sorter100|12982_  = \new_Sorter100|12881_  | \new_Sorter100|12882_ ;
  assign \new_Sorter100|12983_  = \new_Sorter100|12883_  & \new_Sorter100|12884_ ;
  assign \new_Sorter100|12984_  = \new_Sorter100|12883_  | \new_Sorter100|12884_ ;
  assign \new_Sorter100|12985_  = \new_Sorter100|12885_  & \new_Sorter100|12886_ ;
  assign \new_Sorter100|12986_  = \new_Sorter100|12885_  | \new_Sorter100|12886_ ;
  assign \new_Sorter100|12987_  = \new_Sorter100|12887_  & \new_Sorter100|12888_ ;
  assign \new_Sorter100|12988_  = \new_Sorter100|12887_  | \new_Sorter100|12888_ ;
  assign \new_Sorter100|12989_  = \new_Sorter100|12889_  & \new_Sorter100|12890_ ;
  assign \new_Sorter100|12990_  = \new_Sorter100|12889_  | \new_Sorter100|12890_ ;
  assign \new_Sorter100|12991_  = \new_Sorter100|12891_  & \new_Sorter100|12892_ ;
  assign \new_Sorter100|12992_  = \new_Sorter100|12891_  | \new_Sorter100|12892_ ;
  assign \new_Sorter100|12993_  = \new_Sorter100|12893_  & \new_Sorter100|12894_ ;
  assign \new_Sorter100|12994_  = \new_Sorter100|12893_  | \new_Sorter100|12894_ ;
  assign \new_Sorter100|12995_  = \new_Sorter100|12895_  & \new_Sorter100|12896_ ;
  assign \new_Sorter100|12996_  = \new_Sorter100|12895_  | \new_Sorter100|12896_ ;
  assign \new_Sorter100|12997_  = \new_Sorter100|12897_  & \new_Sorter100|12898_ ;
  assign \new_Sorter100|12998_  = \new_Sorter100|12897_  | \new_Sorter100|12898_ ;
  assign \new_Sorter100|13000_  = \new_Sorter100|12900_  & \new_Sorter100|12901_ ;
  assign \new_Sorter100|13001_  = \new_Sorter100|12900_  | \new_Sorter100|12901_ ;
  assign \new_Sorter100|13002_  = \new_Sorter100|12902_  & \new_Sorter100|12903_ ;
  assign \new_Sorter100|13003_  = \new_Sorter100|12902_  | \new_Sorter100|12903_ ;
  assign \new_Sorter100|13004_  = \new_Sorter100|12904_  & \new_Sorter100|12905_ ;
  assign \new_Sorter100|13005_  = \new_Sorter100|12904_  | \new_Sorter100|12905_ ;
  assign \new_Sorter100|13006_  = \new_Sorter100|12906_  & \new_Sorter100|12907_ ;
  assign \new_Sorter100|13007_  = \new_Sorter100|12906_  | \new_Sorter100|12907_ ;
  assign \new_Sorter100|13008_  = \new_Sorter100|12908_  & \new_Sorter100|12909_ ;
  assign \new_Sorter100|13009_  = \new_Sorter100|12908_  | \new_Sorter100|12909_ ;
  assign \new_Sorter100|13010_  = \new_Sorter100|12910_  & \new_Sorter100|12911_ ;
  assign \new_Sorter100|13011_  = \new_Sorter100|12910_  | \new_Sorter100|12911_ ;
  assign \new_Sorter100|13012_  = \new_Sorter100|12912_  & \new_Sorter100|12913_ ;
  assign \new_Sorter100|13013_  = \new_Sorter100|12912_  | \new_Sorter100|12913_ ;
  assign \new_Sorter100|13014_  = \new_Sorter100|12914_  & \new_Sorter100|12915_ ;
  assign \new_Sorter100|13015_  = \new_Sorter100|12914_  | \new_Sorter100|12915_ ;
  assign \new_Sorter100|13016_  = \new_Sorter100|12916_  & \new_Sorter100|12917_ ;
  assign \new_Sorter100|13017_  = \new_Sorter100|12916_  | \new_Sorter100|12917_ ;
  assign \new_Sorter100|13018_  = \new_Sorter100|12918_  & \new_Sorter100|12919_ ;
  assign \new_Sorter100|13019_  = \new_Sorter100|12918_  | \new_Sorter100|12919_ ;
  assign \new_Sorter100|13020_  = \new_Sorter100|12920_  & \new_Sorter100|12921_ ;
  assign \new_Sorter100|13021_  = \new_Sorter100|12920_  | \new_Sorter100|12921_ ;
  assign \new_Sorter100|13022_  = \new_Sorter100|12922_  & \new_Sorter100|12923_ ;
  assign \new_Sorter100|13023_  = \new_Sorter100|12922_  | \new_Sorter100|12923_ ;
  assign \new_Sorter100|13024_  = \new_Sorter100|12924_  & \new_Sorter100|12925_ ;
  assign \new_Sorter100|13025_  = \new_Sorter100|12924_  | \new_Sorter100|12925_ ;
  assign \new_Sorter100|13026_  = \new_Sorter100|12926_  & \new_Sorter100|12927_ ;
  assign \new_Sorter100|13027_  = \new_Sorter100|12926_  | \new_Sorter100|12927_ ;
  assign \new_Sorter100|13028_  = \new_Sorter100|12928_  & \new_Sorter100|12929_ ;
  assign \new_Sorter100|13029_  = \new_Sorter100|12928_  | \new_Sorter100|12929_ ;
  assign \new_Sorter100|13030_  = \new_Sorter100|12930_  & \new_Sorter100|12931_ ;
  assign \new_Sorter100|13031_  = \new_Sorter100|12930_  | \new_Sorter100|12931_ ;
  assign \new_Sorter100|13032_  = \new_Sorter100|12932_  & \new_Sorter100|12933_ ;
  assign \new_Sorter100|13033_  = \new_Sorter100|12932_  | \new_Sorter100|12933_ ;
  assign \new_Sorter100|13034_  = \new_Sorter100|12934_  & \new_Sorter100|12935_ ;
  assign \new_Sorter100|13035_  = \new_Sorter100|12934_  | \new_Sorter100|12935_ ;
  assign \new_Sorter100|13036_  = \new_Sorter100|12936_  & \new_Sorter100|12937_ ;
  assign \new_Sorter100|13037_  = \new_Sorter100|12936_  | \new_Sorter100|12937_ ;
  assign \new_Sorter100|13038_  = \new_Sorter100|12938_  & \new_Sorter100|12939_ ;
  assign \new_Sorter100|13039_  = \new_Sorter100|12938_  | \new_Sorter100|12939_ ;
  assign \new_Sorter100|13040_  = \new_Sorter100|12940_  & \new_Sorter100|12941_ ;
  assign \new_Sorter100|13041_  = \new_Sorter100|12940_  | \new_Sorter100|12941_ ;
  assign \new_Sorter100|13042_  = \new_Sorter100|12942_  & \new_Sorter100|12943_ ;
  assign \new_Sorter100|13043_  = \new_Sorter100|12942_  | \new_Sorter100|12943_ ;
  assign \new_Sorter100|13044_  = \new_Sorter100|12944_  & \new_Sorter100|12945_ ;
  assign \new_Sorter100|13045_  = \new_Sorter100|12944_  | \new_Sorter100|12945_ ;
  assign \new_Sorter100|13046_  = \new_Sorter100|12946_  & \new_Sorter100|12947_ ;
  assign \new_Sorter100|13047_  = \new_Sorter100|12946_  | \new_Sorter100|12947_ ;
  assign \new_Sorter100|13048_  = \new_Sorter100|12948_  & \new_Sorter100|12949_ ;
  assign \new_Sorter100|13049_  = \new_Sorter100|12948_  | \new_Sorter100|12949_ ;
  assign \new_Sorter100|13050_  = \new_Sorter100|12950_  & \new_Sorter100|12951_ ;
  assign \new_Sorter100|13051_  = \new_Sorter100|12950_  | \new_Sorter100|12951_ ;
  assign \new_Sorter100|13052_  = \new_Sorter100|12952_  & \new_Sorter100|12953_ ;
  assign \new_Sorter100|13053_  = \new_Sorter100|12952_  | \new_Sorter100|12953_ ;
  assign \new_Sorter100|13054_  = \new_Sorter100|12954_  & \new_Sorter100|12955_ ;
  assign \new_Sorter100|13055_  = \new_Sorter100|12954_  | \new_Sorter100|12955_ ;
  assign \new_Sorter100|13056_  = \new_Sorter100|12956_  & \new_Sorter100|12957_ ;
  assign \new_Sorter100|13057_  = \new_Sorter100|12956_  | \new_Sorter100|12957_ ;
  assign \new_Sorter100|13058_  = \new_Sorter100|12958_  & \new_Sorter100|12959_ ;
  assign \new_Sorter100|13059_  = \new_Sorter100|12958_  | \new_Sorter100|12959_ ;
  assign \new_Sorter100|13060_  = \new_Sorter100|12960_  & \new_Sorter100|12961_ ;
  assign \new_Sorter100|13061_  = \new_Sorter100|12960_  | \new_Sorter100|12961_ ;
  assign \new_Sorter100|13062_  = \new_Sorter100|12962_  & \new_Sorter100|12963_ ;
  assign \new_Sorter100|13063_  = \new_Sorter100|12962_  | \new_Sorter100|12963_ ;
  assign \new_Sorter100|13064_  = \new_Sorter100|12964_  & \new_Sorter100|12965_ ;
  assign \new_Sorter100|13065_  = \new_Sorter100|12964_  | \new_Sorter100|12965_ ;
  assign \new_Sorter100|13066_  = \new_Sorter100|12966_  & \new_Sorter100|12967_ ;
  assign \new_Sorter100|13067_  = \new_Sorter100|12966_  | \new_Sorter100|12967_ ;
  assign \new_Sorter100|13068_  = \new_Sorter100|12968_  & \new_Sorter100|12969_ ;
  assign \new_Sorter100|13069_  = \new_Sorter100|12968_  | \new_Sorter100|12969_ ;
  assign \new_Sorter100|13070_  = \new_Sorter100|12970_  & \new_Sorter100|12971_ ;
  assign \new_Sorter100|13071_  = \new_Sorter100|12970_  | \new_Sorter100|12971_ ;
  assign \new_Sorter100|13072_  = \new_Sorter100|12972_  & \new_Sorter100|12973_ ;
  assign \new_Sorter100|13073_  = \new_Sorter100|12972_  | \new_Sorter100|12973_ ;
  assign \new_Sorter100|13074_  = \new_Sorter100|12974_  & \new_Sorter100|12975_ ;
  assign \new_Sorter100|13075_  = \new_Sorter100|12974_  | \new_Sorter100|12975_ ;
  assign \new_Sorter100|13076_  = \new_Sorter100|12976_  & \new_Sorter100|12977_ ;
  assign \new_Sorter100|13077_  = \new_Sorter100|12976_  | \new_Sorter100|12977_ ;
  assign \new_Sorter100|13078_  = \new_Sorter100|12978_  & \new_Sorter100|12979_ ;
  assign \new_Sorter100|13079_  = \new_Sorter100|12978_  | \new_Sorter100|12979_ ;
  assign \new_Sorter100|13080_  = \new_Sorter100|12980_  & \new_Sorter100|12981_ ;
  assign \new_Sorter100|13081_  = \new_Sorter100|12980_  | \new_Sorter100|12981_ ;
  assign \new_Sorter100|13082_  = \new_Sorter100|12982_  & \new_Sorter100|12983_ ;
  assign \new_Sorter100|13083_  = \new_Sorter100|12982_  | \new_Sorter100|12983_ ;
  assign \new_Sorter100|13084_  = \new_Sorter100|12984_  & \new_Sorter100|12985_ ;
  assign \new_Sorter100|13085_  = \new_Sorter100|12984_  | \new_Sorter100|12985_ ;
  assign \new_Sorter100|13086_  = \new_Sorter100|12986_  & \new_Sorter100|12987_ ;
  assign \new_Sorter100|13087_  = \new_Sorter100|12986_  | \new_Sorter100|12987_ ;
  assign \new_Sorter100|13088_  = \new_Sorter100|12988_  & \new_Sorter100|12989_ ;
  assign \new_Sorter100|13089_  = \new_Sorter100|12988_  | \new_Sorter100|12989_ ;
  assign \new_Sorter100|13090_  = \new_Sorter100|12990_  & \new_Sorter100|12991_ ;
  assign \new_Sorter100|13091_  = \new_Sorter100|12990_  | \new_Sorter100|12991_ ;
  assign \new_Sorter100|13092_  = \new_Sorter100|12992_  & \new_Sorter100|12993_ ;
  assign \new_Sorter100|13093_  = \new_Sorter100|12992_  | \new_Sorter100|12993_ ;
  assign \new_Sorter100|13094_  = \new_Sorter100|12994_  & \new_Sorter100|12995_ ;
  assign \new_Sorter100|13095_  = \new_Sorter100|12994_  | \new_Sorter100|12995_ ;
  assign \new_Sorter100|13096_  = \new_Sorter100|12996_  & \new_Sorter100|12997_ ;
  assign \new_Sorter100|13097_  = \new_Sorter100|12996_  | \new_Sorter100|12997_ ;
  assign \new_Sorter100|13098_  = \new_Sorter100|12998_  & \new_Sorter100|12999_ ;
  assign \new_Sorter100|13099_  = \new_Sorter100|12998_  | \new_Sorter100|12999_ ;
  assign \new_Sorter100|13100_  = \new_Sorter100|13000_ ;
  assign \new_Sorter100|13199_  = \new_Sorter100|13099_ ;
  assign \new_Sorter100|13101_  = \new_Sorter100|13001_  & \new_Sorter100|13002_ ;
  assign \new_Sorter100|13102_  = \new_Sorter100|13001_  | \new_Sorter100|13002_ ;
  assign \new_Sorter100|13103_  = \new_Sorter100|13003_  & \new_Sorter100|13004_ ;
  assign \new_Sorter100|13104_  = \new_Sorter100|13003_  | \new_Sorter100|13004_ ;
  assign \new_Sorter100|13105_  = \new_Sorter100|13005_  & \new_Sorter100|13006_ ;
  assign \new_Sorter100|13106_  = \new_Sorter100|13005_  | \new_Sorter100|13006_ ;
  assign \new_Sorter100|13107_  = \new_Sorter100|13007_  & \new_Sorter100|13008_ ;
  assign \new_Sorter100|13108_  = \new_Sorter100|13007_  | \new_Sorter100|13008_ ;
  assign \new_Sorter100|13109_  = \new_Sorter100|13009_  & \new_Sorter100|13010_ ;
  assign \new_Sorter100|13110_  = \new_Sorter100|13009_  | \new_Sorter100|13010_ ;
  assign \new_Sorter100|13111_  = \new_Sorter100|13011_  & \new_Sorter100|13012_ ;
  assign \new_Sorter100|13112_  = \new_Sorter100|13011_  | \new_Sorter100|13012_ ;
  assign \new_Sorter100|13113_  = \new_Sorter100|13013_  & \new_Sorter100|13014_ ;
  assign \new_Sorter100|13114_  = \new_Sorter100|13013_  | \new_Sorter100|13014_ ;
  assign \new_Sorter100|13115_  = \new_Sorter100|13015_  & \new_Sorter100|13016_ ;
  assign \new_Sorter100|13116_  = \new_Sorter100|13015_  | \new_Sorter100|13016_ ;
  assign \new_Sorter100|13117_  = \new_Sorter100|13017_  & \new_Sorter100|13018_ ;
  assign \new_Sorter100|13118_  = \new_Sorter100|13017_  | \new_Sorter100|13018_ ;
  assign \new_Sorter100|13119_  = \new_Sorter100|13019_  & \new_Sorter100|13020_ ;
  assign \new_Sorter100|13120_  = \new_Sorter100|13019_  | \new_Sorter100|13020_ ;
  assign \new_Sorter100|13121_  = \new_Sorter100|13021_  & \new_Sorter100|13022_ ;
  assign \new_Sorter100|13122_  = \new_Sorter100|13021_  | \new_Sorter100|13022_ ;
  assign \new_Sorter100|13123_  = \new_Sorter100|13023_  & \new_Sorter100|13024_ ;
  assign \new_Sorter100|13124_  = \new_Sorter100|13023_  | \new_Sorter100|13024_ ;
  assign \new_Sorter100|13125_  = \new_Sorter100|13025_  & \new_Sorter100|13026_ ;
  assign \new_Sorter100|13126_  = \new_Sorter100|13025_  | \new_Sorter100|13026_ ;
  assign \new_Sorter100|13127_  = \new_Sorter100|13027_  & \new_Sorter100|13028_ ;
  assign \new_Sorter100|13128_  = \new_Sorter100|13027_  | \new_Sorter100|13028_ ;
  assign \new_Sorter100|13129_  = \new_Sorter100|13029_  & \new_Sorter100|13030_ ;
  assign \new_Sorter100|13130_  = \new_Sorter100|13029_  | \new_Sorter100|13030_ ;
  assign \new_Sorter100|13131_  = \new_Sorter100|13031_  & \new_Sorter100|13032_ ;
  assign \new_Sorter100|13132_  = \new_Sorter100|13031_  | \new_Sorter100|13032_ ;
  assign \new_Sorter100|13133_  = \new_Sorter100|13033_  & \new_Sorter100|13034_ ;
  assign \new_Sorter100|13134_  = \new_Sorter100|13033_  | \new_Sorter100|13034_ ;
  assign \new_Sorter100|13135_  = \new_Sorter100|13035_  & \new_Sorter100|13036_ ;
  assign \new_Sorter100|13136_  = \new_Sorter100|13035_  | \new_Sorter100|13036_ ;
  assign \new_Sorter100|13137_  = \new_Sorter100|13037_  & \new_Sorter100|13038_ ;
  assign \new_Sorter100|13138_  = \new_Sorter100|13037_  | \new_Sorter100|13038_ ;
  assign \new_Sorter100|13139_  = \new_Sorter100|13039_  & \new_Sorter100|13040_ ;
  assign \new_Sorter100|13140_  = \new_Sorter100|13039_  | \new_Sorter100|13040_ ;
  assign \new_Sorter100|13141_  = \new_Sorter100|13041_  & \new_Sorter100|13042_ ;
  assign \new_Sorter100|13142_  = \new_Sorter100|13041_  | \new_Sorter100|13042_ ;
  assign \new_Sorter100|13143_  = \new_Sorter100|13043_  & \new_Sorter100|13044_ ;
  assign \new_Sorter100|13144_  = \new_Sorter100|13043_  | \new_Sorter100|13044_ ;
  assign \new_Sorter100|13145_  = \new_Sorter100|13045_  & \new_Sorter100|13046_ ;
  assign \new_Sorter100|13146_  = \new_Sorter100|13045_  | \new_Sorter100|13046_ ;
  assign \new_Sorter100|13147_  = \new_Sorter100|13047_  & \new_Sorter100|13048_ ;
  assign \new_Sorter100|13148_  = \new_Sorter100|13047_  | \new_Sorter100|13048_ ;
  assign \new_Sorter100|13149_  = \new_Sorter100|13049_  & \new_Sorter100|13050_ ;
  assign \new_Sorter100|13150_  = \new_Sorter100|13049_  | \new_Sorter100|13050_ ;
  assign \new_Sorter100|13151_  = \new_Sorter100|13051_  & \new_Sorter100|13052_ ;
  assign \new_Sorter100|13152_  = \new_Sorter100|13051_  | \new_Sorter100|13052_ ;
  assign \new_Sorter100|13153_  = \new_Sorter100|13053_  & \new_Sorter100|13054_ ;
  assign \new_Sorter100|13154_  = \new_Sorter100|13053_  | \new_Sorter100|13054_ ;
  assign \new_Sorter100|13155_  = \new_Sorter100|13055_  & \new_Sorter100|13056_ ;
  assign \new_Sorter100|13156_  = \new_Sorter100|13055_  | \new_Sorter100|13056_ ;
  assign \new_Sorter100|13157_  = \new_Sorter100|13057_  & \new_Sorter100|13058_ ;
  assign \new_Sorter100|13158_  = \new_Sorter100|13057_  | \new_Sorter100|13058_ ;
  assign \new_Sorter100|13159_  = \new_Sorter100|13059_  & \new_Sorter100|13060_ ;
  assign \new_Sorter100|13160_  = \new_Sorter100|13059_  | \new_Sorter100|13060_ ;
  assign \new_Sorter100|13161_  = \new_Sorter100|13061_  & \new_Sorter100|13062_ ;
  assign \new_Sorter100|13162_  = \new_Sorter100|13061_  | \new_Sorter100|13062_ ;
  assign \new_Sorter100|13163_  = \new_Sorter100|13063_  & \new_Sorter100|13064_ ;
  assign \new_Sorter100|13164_  = \new_Sorter100|13063_  | \new_Sorter100|13064_ ;
  assign \new_Sorter100|13165_  = \new_Sorter100|13065_  & \new_Sorter100|13066_ ;
  assign \new_Sorter100|13166_  = \new_Sorter100|13065_  | \new_Sorter100|13066_ ;
  assign \new_Sorter100|13167_  = \new_Sorter100|13067_  & \new_Sorter100|13068_ ;
  assign \new_Sorter100|13168_  = \new_Sorter100|13067_  | \new_Sorter100|13068_ ;
  assign \new_Sorter100|13169_  = \new_Sorter100|13069_  & \new_Sorter100|13070_ ;
  assign \new_Sorter100|13170_  = \new_Sorter100|13069_  | \new_Sorter100|13070_ ;
  assign \new_Sorter100|13171_  = \new_Sorter100|13071_  & \new_Sorter100|13072_ ;
  assign \new_Sorter100|13172_  = \new_Sorter100|13071_  | \new_Sorter100|13072_ ;
  assign \new_Sorter100|13173_  = \new_Sorter100|13073_  & \new_Sorter100|13074_ ;
  assign \new_Sorter100|13174_  = \new_Sorter100|13073_  | \new_Sorter100|13074_ ;
  assign \new_Sorter100|13175_  = \new_Sorter100|13075_  & \new_Sorter100|13076_ ;
  assign \new_Sorter100|13176_  = \new_Sorter100|13075_  | \new_Sorter100|13076_ ;
  assign \new_Sorter100|13177_  = \new_Sorter100|13077_  & \new_Sorter100|13078_ ;
  assign \new_Sorter100|13178_  = \new_Sorter100|13077_  | \new_Sorter100|13078_ ;
  assign \new_Sorter100|13179_  = \new_Sorter100|13079_  & \new_Sorter100|13080_ ;
  assign \new_Sorter100|13180_  = \new_Sorter100|13079_  | \new_Sorter100|13080_ ;
  assign \new_Sorter100|13181_  = \new_Sorter100|13081_  & \new_Sorter100|13082_ ;
  assign \new_Sorter100|13182_  = \new_Sorter100|13081_  | \new_Sorter100|13082_ ;
  assign \new_Sorter100|13183_  = \new_Sorter100|13083_  & \new_Sorter100|13084_ ;
  assign \new_Sorter100|13184_  = \new_Sorter100|13083_  | \new_Sorter100|13084_ ;
  assign \new_Sorter100|13185_  = \new_Sorter100|13085_  & \new_Sorter100|13086_ ;
  assign \new_Sorter100|13186_  = \new_Sorter100|13085_  | \new_Sorter100|13086_ ;
  assign \new_Sorter100|13187_  = \new_Sorter100|13087_  & \new_Sorter100|13088_ ;
  assign \new_Sorter100|13188_  = \new_Sorter100|13087_  | \new_Sorter100|13088_ ;
  assign \new_Sorter100|13189_  = \new_Sorter100|13089_  & \new_Sorter100|13090_ ;
  assign \new_Sorter100|13190_  = \new_Sorter100|13089_  | \new_Sorter100|13090_ ;
  assign \new_Sorter100|13191_  = \new_Sorter100|13091_  & \new_Sorter100|13092_ ;
  assign \new_Sorter100|13192_  = \new_Sorter100|13091_  | \new_Sorter100|13092_ ;
  assign \new_Sorter100|13193_  = \new_Sorter100|13093_  & \new_Sorter100|13094_ ;
  assign \new_Sorter100|13194_  = \new_Sorter100|13093_  | \new_Sorter100|13094_ ;
  assign \new_Sorter100|13195_  = \new_Sorter100|13095_  & \new_Sorter100|13096_ ;
  assign \new_Sorter100|13196_  = \new_Sorter100|13095_  | \new_Sorter100|13096_ ;
  assign \new_Sorter100|13197_  = \new_Sorter100|13097_  & \new_Sorter100|13098_ ;
  assign \new_Sorter100|13198_  = \new_Sorter100|13097_  | \new_Sorter100|13098_ ;
  assign \new_Sorter100|13200_  = \new_Sorter100|13100_  & \new_Sorter100|13101_ ;
  assign \new_Sorter100|13201_  = \new_Sorter100|13100_  | \new_Sorter100|13101_ ;
  assign \new_Sorter100|13202_  = \new_Sorter100|13102_  & \new_Sorter100|13103_ ;
  assign \new_Sorter100|13203_  = \new_Sorter100|13102_  | \new_Sorter100|13103_ ;
  assign \new_Sorter100|13204_  = \new_Sorter100|13104_  & \new_Sorter100|13105_ ;
  assign \new_Sorter100|13205_  = \new_Sorter100|13104_  | \new_Sorter100|13105_ ;
  assign \new_Sorter100|13206_  = \new_Sorter100|13106_  & \new_Sorter100|13107_ ;
  assign \new_Sorter100|13207_  = \new_Sorter100|13106_  | \new_Sorter100|13107_ ;
  assign \new_Sorter100|13208_  = \new_Sorter100|13108_  & \new_Sorter100|13109_ ;
  assign \new_Sorter100|13209_  = \new_Sorter100|13108_  | \new_Sorter100|13109_ ;
  assign \new_Sorter100|13210_  = \new_Sorter100|13110_  & \new_Sorter100|13111_ ;
  assign \new_Sorter100|13211_  = \new_Sorter100|13110_  | \new_Sorter100|13111_ ;
  assign \new_Sorter100|13212_  = \new_Sorter100|13112_  & \new_Sorter100|13113_ ;
  assign \new_Sorter100|13213_  = \new_Sorter100|13112_  | \new_Sorter100|13113_ ;
  assign \new_Sorter100|13214_  = \new_Sorter100|13114_  & \new_Sorter100|13115_ ;
  assign \new_Sorter100|13215_  = \new_Sorter100|13114_  | \new_Sorter100|13115_ ;
  assign \new_Sorter100|13216_  = \new_Sorter100|13116_  & \new_Sorter100|13117_ ;
  assign \new_Sorter100|13217_  = \new_Sorter100|13116_  | \new_Sorter100|13117_ ;
  assign \new_Sorter100|13218_  = \new_Sorter100|13118_  & \new_Sorter100|13119_ ;
  assign \new_Sorter100|13219_  = \new_Sorter100|13118_  | \new_Sorter100|13119_ ;
  assign \new_Sorter100|13220_  = \new_Sorter100|13120_  & \new_Sorter100|13121_ ;
  assign \new_Sorter100|13221_  = \new_Sorter100|13120_  | \new_Sorter100|13121_ ;
  assign \new_Sorter100|13222_  = \new_Sorter100|13122_  & \new_Sorter100|13123_ ;
  assign \new_Sorter100|13223_  = \new_Sorter100|13122_  | \new_Sorter100|13123_ ;
  assign \new_Sorter100|13224_  = \new_Sorter100|13124_  & \new_Sorter100|13125_ ;
  assign \new_Sorter100|13225_  = \new_Sorter100|13124_  | \new_Sorter100|13125_ ;
  assign \new_Sorter100|13226_  = \new_Sorter100|13126_  & \new_Sorter100|13127_ ;
  assign \new_Sorter100|13227_  = \new_Sorter100|13126_  | \new_Sorter100|13127_ ;
  assign \new_Sorter100|13228_  = \new_Sorter100|13128_  & \new_Sorter100|13129_ ;
  assign \new_Sorter100|13229_  = \new_Sorter100|13128_  | \new_Sorter100|13129_ ;
  assign \new_Sorter100|13230_  = \new_Sorter100|13130_  & \new_Sorter100|13131_ ;
  assign \new_Sorter100|13231_  = \new_Sorter100|13130_  | \new_Sorter100|13131_ ;
  assign \new_Sorter100|13232_  = \new_Sorter100|13132_  & \new_Sorter100|13133_ ;
  assign \new_Sorter100|13233_  = \new_Sorter100|13132_  | \new_Sorter100|13133_ ;
  assign \new_Sorter100|13234_  = \new_Sorter100|13134_  & \new_Sorter100|13135_ ;
  assign \new_Sorter100|13235_  = \new_Sorter100|13134_  | \new_Sorter100|13135_ ;
  assign \new_Sorter100|13236_  = \new_Sorter100|13136_  & \new_Sorter100|13137_ ;
  assign \new_Sorter100|13237_  = \new_Sorter100|13136_  | \new_Sorter100|13137_ ;
  assign \new_Sorter100|13238_  = \new_Sorter100|13138_  & \new_Sorter100|13139_ ;
  assign \new_Sorter100|13239_  = \new_Sorter100|13138_  | \new_Sorter100|13139_ ;
  assign \new_Sorter100|13240_  = \new_Sorter100|13140_  & \new_Sorter100|13141_ ;
  assign \new_Sorter100|13241_  = \new_Sorter100|13140_  | \new_Sorter100|13141_ ;
  assign \new_Sorter100|13242_  = \new_Sorter100|13142_  & \new_Sorter100|13143_ ;
  assign \new_Sorter100|13243_  = \new_Sorter100|13142_  | \new_Sorter100|13143_ ;
  assign \new_Sorter100|13244_  = \new_Sorter100|13144_  & \new_Sorter100|13145_ ;
  assign \new_Sorter100|13245_  = \new_Sorter100|13144_  | \new_Sorter100|13145_ ;
  assign \new_Sorter100|13246_  = \new_Sorter100|13146_  & \new_Sorter100|13147_ ;
  assign \new_Sorter100|13247_  = \new_Sorter100|13146_  | \new_Sorter100|13147_ ;
  assign \new_Sorter100|13248_  = \new_Sorter100|13148_  & \new_Sorter100|13149_ ;
  assign \new_Sorter100|13249_  = \new_Sorter100|13148_  | \new_Sorter100|13149_ ;
  assign \new_Sorter100|13250_  = \new_Sorter100|13150_  & \new_Sorter100|13151_ ;
  assign \new_Sorter100|13251_  = \new_Sorter100|13150_  | \new_Sorter100|13151_ ;
  assign \new_Sorter100|13252_  = \new_Sorter100|13152_  & \new_Sorter100|13153_ ;
  assign \new_Sorter100|13253_  = \new_Sorter100|13152_  | \new_Sorter100|13153_ ;
  assign \new_Sorter100|13254_  = \new_Sorter100|13154_  & \new_Sorter100|13155_ ;
  assign \new_Sorter100|13255_  = \new_Sorter100|13154_  | \new_Sorter100|13155_ ;
  assign \new_Sorter100|13256_  = \new_Sorter100|13156_  & \new_Sorter100|13157_ ;
  assign \new_Sorter100|13257_  = \new_Sorter100|13156_  | \new_Sorter100|13157_ ;
  assign \new_Sorter100|13258_  = \new_Sorter100|13158_  & \new_Sorter100|13159_ ;
  assign \new_Sorter100|13259_  = \new_Sorter100|13158_  | \new_Sorter100|13159_ ;
  assign \new_Sorter100|13260_  = \new_Sorter100|13160_  & \new_Sorter100|13161_ ;
  assign \new_Sorter100|13261_  = \new_Sorter100|13160_  | \new_Sorter100|13161_ ;
  assign \new_Sorter100|13262_  = \new_Sorter100|13162_  & \new_Sorter100|13163_ ;
  assign \new_Sorter100|13263_  = \new_Sorter100|13162_  | \new_Sorter100|13163_ ;
  assign \new_Sorter100|13264_  = \new_Sorter100|13164_  & \new_Sorter100|13165_ ;
  assign \new_Sorter100|13265_  = \new_Sorter100|13164_  | \new_Sorter100|13165_ ;
  assign \new_Sorter100|13266_  = \new_Sorter100|13166_  & \new_Sorter100|13167_ ;
  assign \new_Sorter100|13267_  = \new_Sorter100|13166_  | \new_Sorter100|13167_ ;
  assign \new_Sorter100|13268_  = \new_Sorter100|13168_  & \new_Sorter100|13169_ ;
  assign \new_Sorter100|13269_  = \new_Sorter100|13168_  | \new_Sorter100|13169_ ;
  assign \new_Sorter100|13270_  = \new_Sorter100|13170_  & \new_Sorter100|13171_ ;
  assign \new_Sorter100|13271_  = \new_Sorter100|13170_  | \new_Sorter100|13171_ ;
  assign \new_Sorter100|13272_  = \new_Sorter100|13172_  & \new_Sorter100|13173_ ;
  assign \new_Sorter100|13273_  = \new_Sorter100|13172_  | \new_Sorter100|13173_ ;
  assign \new_Sorter100|13274_  = \new_Sorter100|13174_  & \new_Sorter100|13175_ ;
  assign \new_Sorter100|13275_  = \new_Sorter100|13174_  | \new_Sorter100|13175_ ;
  assign \new_Sorter100|13276_  = \new_Sorter100|13176_  & \new_Sorter100|13177_ ;
  assign \new_Sorter100|13277_  = \new_Sorter100|13176_  | \new_Sorter100|13177_ ;
  assign \new_Sorter100|13278_  = \new_Sorter100|13178_  & \new_Sorter100|13179_ ;
  assign \new_Sorter100|13279_  = \new_Sorter100|13178_  | \new_Sorter100|13179_ ;
  assign \new_Sorter100|13280_  = \new_Sorter100|13180_  & \new_Sorter100|13181_ ;
  assign \new_Sorter100|13281_  = \new_Sorter100|13180_  | \new_Sorter100|13181_ ;
  assign \new_Sorter100|13282_  = \new_Sorter100|13182_  & \new_Sorter100|13183_ ;
  assign \new_Sorter100|13283_  = \new_Sorter100|13182_  | \new_Sorter100|13183_ ;
  assign \new_Sorter100|13284_  = \new_Sorter100|13184_  & \new_Sorter100|13185_ ;
  assign \new_Sorter100|13285_  = \new_Sorter100|13184_  | \new_Sorter100|13185_ ;
  assign \new_Sorter100|13286_  = \new_Sorter100|13186_  & \new_Sorter100|13187_ ;
  assign \new_Sorter100|13287_  = \new_Sorter100|13186_  | \new_Sorter100|13187_ ;
  assign \new_Sorter100|13288_  = \new_Sorter100|13188_  & \new_Sorter100|13189_ ;
  assign \new_Sorter100|13289_  = \new_Sorter100|13188_  | \new_Sorter100|13189_ ;
  assign \new_Sorter100|13290_  = \new_Sorter100|13190_  & \new_Sorter100|13191_ ;
  assign \new_Sorter100|13291_  = \new_Sorter100|13190_  | \new_Sorter100|13191_ ;
  assign \new_Sorter100|13292_  = \new_Sorter100|13192_  & \new_Sorter100|13193_ ;
  assign \new_Sorter100|13293_  = \new_Sorter100|13192_  | \new_Sorter100|13193_ ;
  assign \new_Sorter100|13294_  = \new_Sorter100|13194_  & \new_Sorter100|13195_ ;
  assign \new_Sorter100|13295_  = \new_Sorter100|13194_  | \new_Sorter100|13195_ ;
  assign \new_Sorter100|13296_  = \new_Sorter100|13196_  & \new_Sorter100|13197_ ;
  assign \new_Sorter100|13297_  = \new_Sorter100|13196_  | \new_Sorter100|13197_ ;
  assign \new_Sorter100|13298_  = \new_Sorter100|13198_  & \new_Sorter100|13199_ ;
  assign \new_Sorter100|13299_  = \new_Sorter100|13198_  | \new_Sorter100|13199_ ;
  assign \new_Sorter100|13300_  = \new_Sorter100|13200_ ;
  assign \new_Sorter100|13399_  = \new_Sorter100|13299_ ;
  assign \new_Sorter100|13301_  = \new_Sorter100|13201_  & \new_Sorter100|13202_ ;
  assign \new_Sorter100|13302_  = \new_Sorter100|13201_  | \new_Sorter100|13202_ ;
  assign \new_Sorter100|13303_  = \new_Sorter100|13203_  & \new_Sorter100|13204_ ;
  assign \new_Sorter100|13304_  = \new_Sorter100|13203_  | \new_Sorter100|13204_ ;
  assign \new_Sorter100|13305_  = \new_Sorter100|13205_  & \new_Sorter100|13206_ ;
  assign \new_Sorter100|13306_  = \new_Sorter100|13205_  | \new_Sorter100|13206_ ;
  assign \new_Sorter100|13307_  = \new_Sorter100|13207_  & \new_Sorter100|13208_ ;
  assign \new_Sorter100|13308_  = \new_Sorter100|13207_  | \new_Sorter100|13208_ ;
  assign \new_Sorter100|13309_  = \new_Sorter100|13209_  & \new_Sorter100|13210_ ;
  assign \new_Sorter100|13310_  = \new_Sorter100|13209_  | \new_Sorter100|13210_ ;
  assign \new_Sorter100|13311_  = \new_Sorter100|13211_  & \new_Sorter100|13212_ ;
  assign \new_Sorter100|13312_  = \new_Sorter100|13211_  | \new_Sorter100|13212_ ;
  assign \new_Sorter100|13313_  = \new_Sorter100|13213_  & \new_Sorter100|13214_ ;
  assign \new_Sorter100|13314_  = \new_Sorter100|13213_  | \new_Sorter100|13214_ ;
  assign \new_Sorter100|13315_  = \new_Sorter100|13215_  & \new_Sorter100|13216_ ;
  assign \new_Sorter100|13316_  = \new_Sorter100|13215_  | \new_Sorter100|13216_ ;
  assign \new_Sorter100|13317_  = \new_Sorter100|13217_  & \new_Sorter100|13218_ ;
  assign \new_Sorter100|13318_  = \new_Sorter100|13217_  | \new_Sorter100|13218_ ;
  assign \new_Sorter100|13319_  = \new_Sorter100|13219_  & \new_Sorter100|13220_ ;
  assign \new_Sorter100|13320_  = \new_Sorter100|13219_  | \new_Sorter100|13220_ ;
  assign \new_Sorter100|13321_  = \new_Sorter100|13221_  & \new_Sorter100|13222_ ;
  assign \new_Sorter100|13322_  = \new_Sorter100|13221_  | \new_Sorter100|13222_ ;
  assign \new_Sorter100|13323_  = \new_Sorter100|13223_  & \new_Sorter100|13224_ ;
  assign \new_Sorter100|13324_  = \new_Sorter100|13223_  | \new_Sorter100|13224_ ;
  assign \new_Sorter100|13325_  = \new_Sorter100|13225_  & \new_Sorter100|13226_ ;
  assign \new_Sorter100|13326_  = \new_Sorter100|13225_  | \new_Sorter100|13226_ ;
  assign \new_Sorter100|13327_  = \new_Sorter100|13227_  & \new_Sorter100|13228_ ;
  assign \new_Sorter100|13328_  = \new_Sorter100|13227_  | \new_Sorter100|13228_ ;
  assign \new_Sorter100|13329_  = \new_Sorter100|13229_  & \new_Sorter100|13230_ ;
  assign \new_Sorter100|13330_  = \new_Sorter100|13229_  | \new_Sorter100|13230_ ;
  assign \new_Sorter100|13331_  = \new_Sorter100|13231_  & \new_Sorter100|13232_ ;
  assign \new_Sorter100|13332_  = \new_Sorter100|13231_  | \new_Sorter100|13232_ ;
  assign \new_Sorter100|13333_  = \new_Sorter100|13233_  & \new_Sorter100|13234_ ;
  assign \new_Sorter100|13334_  = \new_Sorter100|13233_  | \new_Sorter100|13234_ ;
  assign \new_Sorter100|13335_  = \new_Sorter100|13235_  & \new_Sorter100|13236_ ;
  assign \new_Sorter100|13336_  = \new_Sorter100|13235_  | \new_Sorter100|13236_ ;
  assign \new_Sorter100|13337_  = \new_Sorter100|13237_  & \new_Sorter100|13238_ ;
  assign \new_Sorter100|13338_  = \new_Sorter100|13237_  | \new_Sorter100|13238_ ;
  assign \new_Sorter100|13339_  = \new_Sorter100|13239_  & \new_Sorter100|13240_ ;
  assign \new_Sorter100|13340_  = \new_Sorter100|13239_  | \new_Sorter100|13240_ ;
  assign \new_Sorter100|13341_  = \new_Sorter100|13241_  & \new_Sorter100|13242_ ;
  assign \new_Sorter100|13342_  = \new_Sorter100|13241_  | \new_Sorter100|13242_ ;
  assign \new_Sorter100|13343_  = \new_Sorter100|13243_  & \new_Sorter100|13244_ ;
  assign \new_Sorter100|13344_  = \new_Sorter100|13243_  | \new_Sorter100|13244_ ;
  assign \new_Sorter100|13345_  = \new_Sorter100|13245_  & \new_Sorter100|13246_ ;
  assign \new_Sorter100|13346_  = \new_Sorter100|13245_  | \new_Sorter100|13246_ ;
  assign \new_Sorter100|13347_  = \new_Sorter100|13247_  & \new_Sorter100|13248_ ;
  assign \new_Sorter100|13348_  = \new_Sorter100|13247_  | \new_Sorter100|13248_ ;
  assign \new_Sorter100|13349_  = \new_Sorter100|13249_  & \new_Sorter100|13250_ ;
  assign \new_Sorter100|13350_  = \new_Sorter100|13249_  | \new_Sorter100|13250_ ;
  assign \new_Sorter100|13351_  = \new_Sorter100|13251_  & \new_Sorter100|13252_ ;
  assign \new_Sorter100|13352_  = \new_Sorter100|13251_  | \new_Sorter100|13252_ ;
  assign \new_Sorter100|13353_  = \new_Sorter100|13253_  & \new_Sorter100|13254_ ;
  assign \new_Sorter100|13354_  = \new_Sorter100|13253_  | \new_Sorter100|13254_ ;
  assign \new_Sorter100|13355_  = \new_Sorter100|13255_  & \new_Sorter100|13256_ ;
  assign \new_Sorter100|13356_  = \new_Sorter100|13255_  | \new_Sorter100|13256_ ;
  assign \new_Sorter100|13357_  = \new_Sorter100|13257_  & \new_Sorter100|13258_ ;
  assign \new_Sorter100|13358_  = \new_Sorter100|13257_  | \new_Sorter100|13258_ ;
  assign \new_Sorter100|13359_  = \new_Sorter100|13259_  & \new_Sorter100|13260_ ;
  assign \new_Sorter100|13360_  = \new_Sorter100|13259_  | \new_Sorter100|13260_ ;
  assign \new_Sorter100|13361_  = \new_Sorter100|13261_  & \new_Sorter100|13262_ ;
  assign \new_Sorter100|13362_  = \new_Sorter100|13261_  | \new_Sorter100|13262_ ;
  assign \new_Sorter100|13363_  = \new_Sorter100|13263_  & \new_Sorter100|13264_ ;
  assign \new_Sorter100|13364_  = \new_Sorter100|13263_  | \new_Sorter100|13264_ ;
  assign \new_Sorter100|13365_  = \new_Sorter100|13265_  & \new_Sorter100|13266_ ;
  assign \new_Sorter100|13366_  = \new_Sorter100|13265_  | \new_Sorter100|13266_ ;
  assign \new_Sorter100|13367_  = \new_Sorter100|13267_  & \new_Sorter100|13268_ ;
  assign \new_Sorter100|13368_  = \new_Sorter100|13267_  | \new_Sorter100|13268_ ;
  assign \new_Sorter100|13369_  = \new_Sorter100|13269_  & \new_Sorter100|13270_ ;
  assign \new_Sorter100|13370_  = \new_Sorter100|13269_  | \new_Sorter100|13270_ ;
  assign \new_Sorter100|13371_  = \new_Sorter100|13271_  & \new_Sorter100|13272_ ;
  assign \new_Sorter100|13372_  = \new_Sorter100|13271_  | \new_Sorter100|13272_ ;
  assign \new_Sorter100|13373_  = \new_Sorter100|13273_  & \new_Sorter100|13274_ ;
  assign \new_Sorter100|13374_  = \new_Sorter100|13273_  | \new_Sorter100|13274_ ;
  assign \new_Sorter100|13375_  = \new_Sorter100|13275_  & \new_Sorter100|13276_ ;
  assign \new_Sorter100|13376_  = \new_Sorter100|13275_  | \new_Sorter100|13276_ ;
  assign \new_Sorter100|13377_  = \new_Sorter100|13277_  & \new_Sorter100|13278_ ;
  assign \new_Sorter100|13378_  = \new_Sorter100|13277_  | \new_Sorter100|13278_ ;
  assign \new_Sorter100|13379_  = \new_Sorter100|13279_  & \new_Sorter100|13280_ ;
  assign \new_Sorter100|13380_  = \new_Sorter100|13279_  | \new_Sorter100|13280_ ;
  assign \new_Sorter100|13381_  = \new_Sorter100|13281_  & \new_Sorter100|13282_ ;
  assign \new_Sorter100|13382_  = \new_Sorter100|13281_  | \new_Sorter100|13282_ ;
  assign \new_Sorter100|13383_  = \new_Sorter100|13283_  & \new_Sorter100|13284_ ;
  assign \new_Sorter100|13384_  = \new_Sorter100|13283_  | \new_Sorter100|13284_ ;
  assign \new_Sorter100|13385_  = \new_Sorter100|13285_  & \new_Sorter100|13286_ ;
  assign \new_Sorter100|13386_  = \new_Sorter100|13285_  | \new_Sorter100|13286_ ;
  assign \new_Sorter100|13387_  = \new_Sorter100|13287_  & \new_Sorter100|13288_ ;
  assign \new_Sorter100|13388_  = \new_Sorter100|13287_  | \new_Sorter100|13288_ ;
  assign \new_Sorter100|13389_  = \new_Sorter100|13289_  & \new_Sorter100|13290_ ;
  assign \new_Sorter100|13390_  = \new_Sorter100|13289_  | \new_Sorter100|13290_ ;
  assign \new_Sorter100|13391_  = \new_Sorter100|13291_  & \new_Sorter100|13292_ ;
  assign \new_Sorter100|13392_  = \new_Sorter100|13291_  | \new_Sorter100|13292_ ;
  assign \new_Sorter100|13393_  = \new_Sorter100|13293_  & \new_Sorter100|13294_ ;
  assign \new_Sorter100|13394_  = \new_Sorter100|13293_  | \new_Sorter100|13294_ ;
  assign \new_Sorter100|13395_  = \new_Sorter100|13295_  & \new_Sorter100|13296_ ;
  assign \new_Sorter100|13396_  = \new_Sorter100|13295_  | \new_Sorter100|13296_ ;
  assign \new_Sorter100|13397_  = \new_Sorter100|13297_  & \new_Sorter100|13298_ ;
  assign \new_Sorter100|13398_  = \new_Sorter100|13297_  | \new_Sorter100|13298_ ;
  assign \new_Sorter100|13400_  = \new_Sorter100|13300_  & \new_Sorter100|13301_ ;
  assign \new_Sorter100|13401_  = \new_Sorter100|13300_  | \new_Sorter100|13301_ ;
  assign \new_Sorter100|13402_  = \new_Sorter100|13302_  & \new_Sorter100|13303_ ;
  assign \new_Sorter100|13403_  = \new_Sorter100|13302_  | \new_Sorter100|13303_ ;
  assign \new_Sorter100|13404_  = \new_Sorter100|13304_  & \new_Sorter100|13305_ ;
  assign \new_Sorter100|13405_  = \new_Sorter100|13304_  | \new_Sorter100|13305_ ;
  assign \new_Sorter100|13406_  = \new_Sorter100|13306_  & \new_Sorter100|13307_ ;
  assign \new_Sorter100|13407_  = \new_Sorter100|13306_  | \new_Sorter100|13307_ ;
  assign \new_Sorter100|13408_  = \new_Sorter100|13308_  & \new_Sorter100|13309_ ;
  assign \new_Sorter100|13409_  = \new_Sorter100|13308_  | \new_Sorter100|13309_ ;
  assign \new_Sorter100|13410_  = \new_Sorter100|13310_  & \new_Sorter100|13311_ ;
  assign \new_Sorter100|13411_  = \new_Sorter100|13310_  | \new_Sorter100|13311_ ;
  assign \new_Sorter100|13412_  = \new_Sorter100|13312_  & \new_Sorter100|13313_ ;
  assign \new_Sorter100|13413_  = \new_Sorter100|13312_  | \new_Sorter100|13313_ ;
  assign \new_Sorter100|13414_  = \new_Sorter100|13314_  & \new_Sorter100|13315_ ;
  assign \new_Sorter100|13415_  = \new_Sorter100|13314_  | \new_Sorter100|13315_ ;
  assign \new_Sorter100|13416_  = \new_Sorter100|13316_  & \new_Sorter100|13317_ ;
  assign \new_Sorter100|13417_  = \new_Sorter100|13316_  | \new_Sorter100|13317_ ;
  assign \new_Sorter100|13418_  = \new_Sorter100|13318_  & \new_Sorter100|13319_ ;
  assign \new_Sorter100|13419_  = \new_Sorter100|13318_  | \new_Sorter100|13319_ ;
  assign \new_Sorter100|13420_  = \new_Sorter100|13320_  & \new_Sorter100|13321_ ;
  assign \new_Sorter100|13421_  = \new_Sorter100|13320_  | \new_Sorter100|13321_ ;
  assign \new_Sorter100|13422_  = \new_Sorter100|13322_  & \new_Sorter100|13323_ ;
  assign \new_Sorter100|13423_  = \new_Sorter100|13322_  | \new_Sorter100|13323_ ;
  assign \new_Sorter100|13424_  = \new_Sorter100|13324_  & \new_Sorter100|13325_ ;
  assign \new_Sorter100|13425_  = \new_Sorter100|13324_  | \new_Sorter100|13325_ ;
  assign \new_Sorter100|13426_  = \new_Sorter100|13326_  & \new_Sorter100|13327_ ;
  assign \new_Sorter100|13427_  = \new_Sorter100|13326_  | \new_Sorter100|13327_ ;
  assign \new_Sorter100|13428_  = \new_Sorter100|13328_  & \new_Sorter100|13329_ ;
  assign \new_Sorter100|13429_  = \new_Sorter100|13328_  | \new_Sorter100|13329_ ;
  assign \new_Sorter100|13430_  = \new_Sorter100|13330_  & \new_Sorter100|13331_ ;
  assign \new_Sorter100|13431_  = \new_Sorter100|13330_  | \new_Sorter100|13331_ ;
  assign \new_Sorter100|13432_  = \new_Sorter100|13332_  & \new_Sorter100|13333_ ;
  assign \new_Sorter100|13433_  = \new_Sorter100|13332_  | \new_Sorter100|13333_ ;
  assign \new_Sorter100|13434_  = \new_Sorter100|13334_  & \new_Sorter100|13335_ ;
  assign \new_Sorter100|13435_  = \new_Sorter100|13334_  | \new_Sorter100|13335_ ;
  assign \new_Sorter100|13436_  = \new_Sorter100|13336_  & \new_Sorter100|13337_ ;
  assign \new_Sorter100|13437_  = \new_Sorter100|13336_  | \new_Sorter100|13337_ ;
  assign \new_Sorter100|13438_  = \new_Sorter100|13338_  & \new_Sorter100|13339_ ;
  assign \new_Sorter100|13439_  = \new_Sorter100|13338_  | \new_Sorter100|13339_ ;
  assign \new_Sorter100|13440_  = \new_Sorter100|13340_  & \new_Sorter100|13341_ ;
  assign \new_Sorter100|13441_  = \new_Sorter100|13340_  | \new_Sorter100|13341_ ;
  assign \new_Sorter100|13442_  = \new_Sorter100|13342_  & \new_Sorter100|13343_ ;
  assign \new_Sorter100|13443_  = \new_Sorter100|13342_  | \new_Sorter100|13343_ ;
  assign \new_Sorter100|13444_  = \new_Sorter100|13344_  & \new_Sorter100|13345_ ;
  assign \new_Sorter100|13445_  = \new_Sorter100|13344_  | \new_Sorter100|13345_ ;
  assign \new_Sorter100|13446_  = \new_Sorter100|13346_  & \new_Sorter100|13347_ ;
  assign \new_Sorter100|13447_  = \new_Sorter100|13346_  | \new_Sorter100|13347_ ;
  assign \new_Sorter100|13448_  = \new_Sorter100|13348_  & \new_Sorter100|13349_ ;
  assign \new_Sorter100|13449_  = \new_Sorter100|13348_  | \new_Sorter100|13349_ ;
  assign \new_Sorter100|13450_  = \new_Sorter100|13350_  & \new_Sorter100|13351_ ;
  assign \new_Sorter100|13451_  = \new_Sorter100|13350_  | \new_Sorter100|13351_ ;
  assign \new_Sorter100|13452_  = \new_Sorter100|13352_  & \new_Sorter100|13353_ ;
  assign \new_Sorter100|13453_  = \new_Sorter100|13352_  | \new_Sorter100|13353_ ;
  assign \new_Sorter100|13454_  = \new_Sorter100|13354_  & \new_Sorter100|13355_ ;
  assign \new_Sorter100|13455_  = \new_Sorter100|13354_  | \new_Sorter100|13355_ ;
  assign \new_Sorter100|13456_  = \new_Sorter100|13356_  & \new_Sorter100|13357_ ;
  assign \new_Sorter100|13457_  = \new_Sorter100|13356_  | \new_Sorter100|13357_ ;
  assign \new_Sorter100|13458_  = \new_Sorter100|13358_  & \new_Sorter100|13359_ ;
  assign \new_Sorter100|13459_  = \new_Sorter100|13358_  | \new_Sorter100|13359_ ;
  assign \new_Sorter100|13460_  = \new_Sorter100|13360_  & \new_Sorter100|13361_ ;
  assign \new_Sorter100|13461_  = \new_Sorter100|13360_  | \new_Sorter100|13361_ ;
  assign \new_Sorter100|13462_  = \new_Sorter100|13362_  & \new_Sorter100|13363_ ;
  assign \new_Sorter100|13463_  = \new_Sorter100|13362_  | \new_Sorter100|13363_ ;
  assign \new_Sorter100|13464_  = \new_Sorter100|13364_  & \new_Sorter100|13365_ ;
  assign \new_Sorter100|13465_  = \new_Sorter100|13364_  | \new_Sorter100|13365_ ;
  assign \new_Sorter100|13466_  = \new_Sorter100|13366_  & \new_Sorter100|13367_ ;
  assign \new_Sorter100|13467_  = \new_Sorter100|13366_  | \new_Sorter100|13367_ ;
  assign \new_Sorter100|13468_  = \new_Sorter100|13368_  & \new_Sorter100|13369_ ;
  assign \new_Sorter100|13469_  = \new_Sorter100|13368_  | \new_Sorter100|13369_ ;
  assign \new_Sorter100|13470_  = \new_Sorter100|13370_  & \new_Sorter100|13371_ ;
  assign \new_Sorter100|13471_  = \new_Sorter100|13370_  | \new_Sorter100|13371_ ;
  assign \new_Sorter100|13472_  = \new_Sorter100|13372_  & \new_Sorter100|13373_ ;
  assign \new_Sorter100|13473_  = \new_Sorter100|13372_  | \new_Sorter100|13373_ ;
  assign \new_Sorter100|13474_  = \new_Sorter100|13374_  & \new_Sorter100|13375_ ;
  assign \new_Sorter100|13475_  = \new_Sorter100|13374_  | \new_Sorter100|13375_ ;
  assign \new_Sorter100|13476_  = \new_Sorter100|13376_  & \new_Sorter100|13377_ ;
  assign \new_Sorter100|13477_  = \new_Sorter100|13376_  | \new_Sorter100|13377_ ;
  assign \new_Sorter100|13478_  = \new_Sorter100|13378_  & \new_Sorter100|13379_ ;
  assign \new_Sorter100|13479_  = \new_Sorter100|13378_  | \new_Sorter100|13379_ ;
  assign \new_Sorter100|13480_  = \new_Sorter100|13380_  & \new_Sorter100|13381_ ;
  assign \new_Sorter100|13481_  = \new_Sorter100|13380_  | \new_Sorter100|13381_ ;
  assign \new_Sorter100|13482_  = \new_Sorter100|13382_  & \new_Sorter100|13383_ ;
  assign \new_Sorter100|13483_  = \new_Sorter100|13382_  | \new_Sorter100|13383_ ;
  assign \new_Sorter100|13484_  = \new_Sorter100|13384_  & \new_Sorter100|13385_ ;
  assign \new_Sorter100|13485_  = \new_Sorter100|13384_  | \new_Sorter100|13385_ ;
  assign \new_Sorter100|13486_  = \new_Sorter100|13386_  & \new_Sorter100|13387_ ;
  assign \new_Sorter100|13487_  = \new_Sorter100|13386_  | \new_Sorter100|13387_ ;
  assign \new_Sorter100|13488_  = \new_Sorter100|13388_  & \new_Sorter100|13389_ ;
  assign \new_Sorter100|13489_  = \new_Sorter100|13388_  | \new_Sorter100|13389_ ;
  assign \new_Sorter100|13490_  = \new_Sorter100|13390_  & \new_Sorter100|13391_ ;
  assign \new_Sorter100|13491_  = \new_Sorter100|13390_  | \new_Sorter100|13391_ ;
  assign \new_Sorter100|13492_  = \new_Sorter100|13392_  & \new_Sorter100|13393_ ;
  assign \new_Sorter100|13493_  = \new_Sorter100|13392_  | \new_Sorter100|13393_ ;
  assign \new_Sorter100|13494_  = \new_Sorter100|13394_  & \new_Sorter100|13395_ ;
  assign \new_Sorter100|13495_  = \new_Sorter100|13394_  | \new_Sorter100|13395_ ;
  assign \new_Sorter100|13496_  = \new_Sorter100|13396_  & \new_Sorter100|13397_ ;
  assign \new_Sorter100|13497_  = \new_Sorter100|13396_  | \new_Sorter100|13397_ ;
  assign \new_Sorter100|13498_  = \new_Sorter100|13398_  & \new_Sorter100|13399_ ;
  assign \new_Sorter100|13499_  = \new_Sorter100|13398_  | \new_Sorter100|13399_ ;
  assign \new_Sorter100|13500_  = \new_Sorter100|13400_ ;
  assign \new_Sorter100|13599_  = \new_Sorter100|13499_ ;
  assign \new_Sorter100|13501_  = \new_Sorter100|13401_  & \new_Sorter100|13402_ ;
  assign \new_Sorter100|13502_  = \new_Sorter100|13401_  | \new_Sorter100|13402_ ;
  assign \new_Sorter100|13503_  = \new_Sorter100|13403_  & \new_Sorter100|13404_ ;
  assign \new_Sorter100|13504_  = \new_Sorter100|13403_  | \new_Sorter100|13404_ ;
  assign \new_Sorter100|13505_  = \new_Sorter100|13405_  & \new_Sorter100|13406_ ;
  assign \new_Sorter100|13506_  = \new_Sorter100|13405_  | \new_Sorter100|13406_ ;
  assign \new_Sorter100|13507_  = \new_Sorter100|13407_  & \new_Sorter100|13408_ ;
  assign \new_Sorter100|13508_  = \new_Sorter100|13407_  | \new_Sorter100|13408_ ;
  assign \new_Sorter100|13509_  = \new_Sorter100|13409_  & \new_Sorter100|13410_ ;
  assign \new_Sorter100|13510_  = \new_Sorter100|13409_  | \new_Sorter100|13410_ ;
  assign \new_Sorter100|13511_  = \new_Sorter100|13411_  & \new_Sorter100|13412_ ;
  assign \new_Sorter100|13512_  = \new_Sorter100|13411_  | \new_Sorter100|13412_ ;
  assign \new_Sorter100|13513_  = \new_Sorter100|13413_  & \new_Sorter100|13414_ ;
  assign \new_Sorter100|13514_  = \new_Sorter100|13413_  | \new_Sorter100|13414_ ;
  assign \new_Sorter100|13515_  = \new_Sorter100|13415_  & \new_Sorter100|13416_ ;
  assign \new_Sorter100|13516_  = \new_Sorter100|13415_  | \new_Sorter100|13416_ ;
  assign \new_Sorter100|13517_  = \new_Sorter100|13417_  & \new_Sorter100|13418_ ;
  assign \new_Sorter100|13518_  = \new_Sorter100|13417_  | \new_Sorter100|13418_ ;
  assign \new_Sorter100|13519_  = \new_Sorter100|13419_  & \new_Sorter100|13420_ ;
  assign \new_Sorter100|13520_  = \new_Sorter100|13419_  | \new_Sorter100|13420_ ;
  assign \new_Sorter100|13521_  = \new_Sorter100|13421_  & \new_Sorter100|13422_ ;
  assign \new_Sorter100|13522_  = \new_Sorter100|13421_  | \new_Sorter100|13422_ ;
  assign \new_Sorter100|13523_  = \new_Sorter100|13423_  & \new_Sorter100|13424_ ;
  assign \new_Sorter100|13524_  = \new_Sorter100|13423_  | \new_Sorter100|13424_ ;
  assign \new_Sorter100|13525_  = \new_Sorter100|13425_  & \new_Sorter100|13426_ ;
  assign \new_Sorter100|13526_  = \new_Sorter100|13425_  | \new_Sorter100|13426_ ;
  assign \new_Sorter100|13527_  = \new_Sorter100|13427_  & \new_Sorter100|13428_ ;
  assign \new_Sorter100|13528_  = \new_Sorter100|13427_  | \new_Sorter100|13428_ ;
  assign \new_Sorter100|13529_  = \new_Sorter100|13429_  & \new_Sorter100|13430_ ;
  assign \new_Sorter100|13530_  = \new_Sorter100|13429_  | \new_Sorter100|13430_ ;
  assign \new_Sorter100|13531_  = \new_Sorter100|13431_  & \new_Sorter100|13432_ ;
  assign \new_Sorter100|13532_  = \new_Sorter100|13431_  | \new_Sorter100|13432_ ;
  assign \new_Sorter100|13533_  = \new_Sorter100|13433_  & \new_Sorter100|13434_ ;
  assign \new_Sorter100|13534_  = \new_Sorter100|13433_  | \new_Sorter100|13434_ ;
  assign \new_Sorter100|13535_  = \new_Sorter100|13435_  & \new_Sorter100|13436_ ;
  assign \new_Sorter100|13536_  = \new_Sorter100|13435_  | \new_Sorter100|13436_ ;
  assign \new_Sorter100|13537_  = \new_Sorter100|13437_  & \new_Sorter100|13438_ ;
  assign \new_Sorter100|13538_  = \new_Sorter100|13437_  | \new_Sorter100|13438_ ;
  assign \new_Sorter100|13539_  = \new_Sorter100|13439_  & \new_Sorter100|13440_ ;
  assign \new_Sorter100|13540_  = \new_Sorter100|13439_  | \new_Sorter100|13440_ ;
  assign \new_Sorter100|13541_  = \new_Sorter100|13441_  & \new_Sorter100|13442_ ;
  assign \new_Sorter100|13542_  = \new_Sorter100|13441_  | \new_Sorter100|13442_ ;
  assign \new_Sorter100|13543_  = \new_Sorter100|13443_  & \new_Sorter100|13444_ ;
  assign \new_Sorter100|13544_  = \new_Sorter100|13443_  | \new_Sorter100|13444_ ;
  assign \new_Sorter100|13545_  = \new_Sorter100|13445_  & \new_Sorter100|13446_ ;
  assign \new_Sorter100|13546_  = \new_Sorter100|13445_  | \new_Sorter100|13446_ ;
  assign \new_Sorter100|13547_  = \new_Sorter100|13447_  & \new_Sorter100|13448_ ;
  assign \new_Sorter100|13548_  = \new_Sorter100|13447_  | \new_Sorter100|13448_ ;
  assign \new_Sorter100|13549_  = \new_Sorter100|13449_  & \new_Sorter100|13450_ ;
  assign \new_Sorter100|13550_  = \new_Sorter100|13449_  | \new_Sorter100|13450_ ;
  assign \new_Sorter100|13551_  = \new_Sorter100|13451_  & \new_Sorter100|13452_ ;
  assign \new_Sorter100|13552_  = \new_Sorter100|13451_  | \new_Sorter100|13452_ ;
  assign \new_Sorter100|13553_  = \new_Sorter100|13453_  & \new_Sorter100|13454_ ;
  assign \new_Sorter100|13554_  = \new_Sorter100|13453_  | \new_Sorter100|13454_ ;
  assign \new_Sorter100|13555_  = \new_Sorter100|13455_  & \new_Sorter100|13456_ ;
  assign \new_Sorter100|13556_  = \new_Sorter100|13455_  | \new_Sorter100|13456_ ;
  assign \new_Sorter100|13557_  = \new_Sorter100|13457_  & \new_Sorter100|13458_ ;
  assign \new_Sorter100|13558_  = \new_Sorter100|13457_  | \new_Sorter100|13458_ ;
  assign \new_Sorter100|13559_  = \new_Sorter100|13459_  & \new_Sorter100|13460_ ;
  assign \new_Sorter100|13560_  = \new_Sorter100|13459_  | \new_Sorter100|13460_ ;
  assign \new_Sorter100|13561_  = \new_Sorter100|13461_  & \new_Sorter100|13462_ ;
  assign \new_Sorter100|13562_  = \new_Sorter100|13461_  | \new_Sorter100|13462_ ;
  assign \new_Sorter100|13563_  = \new_Sorter100|13463_  & \new_Sorter100|13464_ ;
  assign \new_Sorter100|13564_  = \new_Sorter100|13463_  | \new_Sorter100|13464_ ;
  assign \new_Sorter100|13565_  = \new_Sorter100|13465_  & \new_Sorter100|13466_ ;
  assign \new_Sorter100|13566_  = \new_Sorter100|13465_  | \new_Sorter100|13466_ ;
  assign \new_Sorter100|13567_  = \new_Sorter100|13467_  & \new_Sorter100|13468_ ;
  assign \new_Sorter100|13568_  = \new_Sorter100|13467_  | \new_Sorter100|13468_ ;
  assign \new_Sorter100|13569_  = \new_Sorter100|13469_  & \new_Sorter100|13470_ ;
  assign \new_Sorter100|13570_  = \new_Sorter100|13469_  | \new_Sorter100|13470_ ;
  assign \new_Sorter100|13571_  = \new_Sorter100|13471_  & \new_Sorter100|13472_ ;
  assign \new_Sorter100|13572_  = \new_Sorter100|13471_  | \new_Sorter100|13472_ ;
  assign \new_Sorter100|13573_  = \new_Sorter100|13473_  & \new_Sorter100|13474_ ;
  assign \new_Sorter100|13574_  = \new_Sorter100|13473_  | \new_Sorter100|13474_ ;
  assign \new_Sorter100|13575_  = \new_Sorter100|13475_  & \new_Sorter100|13476_ ;
  assign \new_Sorter100|13576_  = \new_Sorter100|13475_  | \new_Sorter100|13476_ ;
  assign \new_Sorter100|13577_  = \new_Sorter100|13477_  & \new_Sorter100|13478_ ;
  assign \new_Sorter100|13578_  = \new_Sorter100|13477_  | \new_Sorter100|13478_ ;
  assign \new_Sorter100|13579_  = \new_Sorter100|13479_  & \new_Sorter100|13480_ ;
  assign \new_Sorter100|13580_  = \new_Sorter100|13479_  | \new_Sorter100|13480_ ;
  assign \new_Sorter100|13581_  = \new_Sorter100|13481_  & \new_Sorter100|13482_ ;
  assign \new_Sorter100|13582_  = \new_Sorter100|13481_  | \new_Sorter100|13482_ ;
  assign \new_Sorter100|13583_  = \new_Sorter100|13483_  & \new_Sorter100|13484_ ;
  assign \new_Sorter100|13584_  = \new_Sorter100|13483_  | \new_Sorter100|13484_ ;
  assign \new_Sorter100|13585_  = \new_Sorter100|13485_  & \new_Sorter100|13486_ ;
  assign \new_Sorter100|13586_  = \new_Sorter100|13485_  | \new_Sorter100|13486_ ;
  assign \new_Sorter100|13587_  = \new_Sorter100|13487_  & \new_Sorter100|13488_ ;
  assign \new_Sorter100|13588_  = \new_Sorter100|13487_  | \new_Sorter100|13488_ ;
  assign \new_Sorter100|13589_  = \new_Sorter100|13489_  & \new_Sorter100|13490_ ;
  assign \new_Sorter100|13590_  = \new_Sorter100|13489_  | \new_Sorter100|13490_ ;
  assign \new_Sorter100|13591_  = \new_Sorter100|13491_  & \new_Sorter100|13492_ ;
  assign \new_Sorter100|13592_  = \new_Sorter100|13491_  | \new_Sorter100|13492_ ;
  assign \new_Sorter100|13593_  = \new_Sorter100|13493_  & \new_Sorter100|13494_ ;
  assign \new_Sorter100|13594_  = \new_Sorter100|13493_  | \new_Sorter100|13494_ ;
  assign \new_Sorter100|13595_  = \new_Sorter100|13495_  & \new_Sorter100|13496_ ;
  assign \new_Sorter100|13596_  = \new_Sorter100|13495_  | \new_Sorter100|13496_ ;
  assign \new_Sorter100|13597_  = \new_Sorter100|13497_  & \new_Sorter100|13498_ ;
  assign \new_Sorter100|13598_  = \new_Sorter100|13497_  | \new_Sorter100|13498_ ;
  assign \new_Sorter100|13600_  = \new_Sorter100|13500_  & \new_Sorter100|13501_ ;
  assign \new_Sorter100|13601_  = \new_Sorter100|13500_  | \new_Sorter100|13501_ ;
  assign \new_Sorter100|13602_  = \new_Sorter100|13502_  & \new_Sorter100|13503_ ;
  assign \new_Sorter100|13603_  = \new_Sorter100|13502_  | \new_Sorter100|13503_ ;
  assign \new_Sorter100|13604_  = \new_Sorter100|13504_  & \new_Sorter100|13505_ ;
  assign \new_Sorter100|13605_  = \new_Sorter100|13504_  | \new_Sorter100|13505_ ;
  assign \new_Sorter100|13606_  = \new_Sorter100|13506_  & \new_Sorter100|13507_ ;
  assign \new_Sorter100|13607_  = \new_Sorter100|13506_  | \new_Sorter100|13507_ ;
  assign \new_Sorter100|13608_  = \new_Sorter100|13508_  & \new_Sorter100|13509_ ;
  assign \new_Sorter100|13609_  = \new_Sorter100|13508_  | \new_Sorter100|13509_ ;
  assign \new_Sorter100|13610_  = \new_Sorter100|13510_  & \new_Sorter100|13511_ ;
  assign \new_Sorter100|13611_  = \new_Sorter100|13510_  | \new_Sorter100|13511_ ;
  assign \new_Sorter100|13612_  = \new_Sorter100|13512_  & \new_Sorter100|13513_ ;
  assign \new_Sorter100|13613_  = \new_Sorter100|13512_  | \new_Sorter100|13513_ ;
  assign \new_Sorter100|13614_  = \new_Sorter100|13514_  & \new_Sorter100|13515_ ;
  assign \new_Sorter100|13615_  = \new_Sorter100|13514_  | \new_Sorter100|13515_ ;
  assign \new_Sorter100|13616_  = \new_Sorter100|13516_  & \new_Sorter100|13517_ ;
  assign \new_Sorter100|13617_  = \new_Sorter100|13516_  | \new_Sorter100|13517_ ;
  assign \new_Sorter100|13618_  = \new_Sorter100|13518_  & \new_Sorter100|13519_ ;
  assign \new_Sorter100|13619_  = \new_Sorter100|13518_  | \new_Sorter100|13519_ ;
  assign \new_Sorter100|13620_  = \new_Sorter100|13520_  & \new_Sorter100|13521_ ;
  assign \new_Sorter100|13621_  = \new_Sorter100|13520_  | \new_Sorter100|13521_ ;
  assign \new_Sorter100|13622_  = \new_Sorter100|13522_  & \new_Sorter100|13523_ ;
  assign \new_Sorter100|13623_  = \new_Sorter100|13522_  | \new_Sorter100|13523_ ;
  assign \new_Sorter100|13624_  = \new_Sorter100|13524_  & \new_Sorter100|13525_ ;
  assign \new_Sorter100|13625_  = \new_Sorter100|13524_  | \new_Sorter100|13525_ ;
  assign \new_Sorter100|13626_  = \new_Sorter100|13526_  & \new_Sorter100|13527_ ;
  assign \new_Sorter100|13627_  = \new_Sorter100|13526_  | \new_Sorter100|13527_ ;
  assign \new_Sorter100|13628_  = \new_Sorter100|13528_  & \new_Sorter100|13529_ ;
  assign \new_Sorter100|13629_  = \new_Sorter100|13528_  | \new_Sorter100|13529_ ;
  assign \new_Sorter100|13630_  = \new_Sorter100|13530_  & \new_Sorter100|13531_ ;
  assign \new_Sorter100|13631_  = \new_Sorter100|13530_  | \new_Sorter100|13531_ ;
  assign \new_Sorter100|13632_  = \new_Sorter100|13532_  & \new_Sorter100|13533_ ;
  assign \new_Sorter100|13633_  = \new_Sorter100|13532_  | \new_Sorter100|13533_ ;
  assign \new_Sorter100|13634_  = \new_Sorter100|13534_  & \new_Sorter100|13535_ ;
  assign \new_Sorter100|13635_  = \new_Sorter100|13534_  | \new_Sorter100|13535_ ;
  assign \new_Sorter100|13636_  = \new_Sorter100|13536_  & \new_Sorter100|13537_ ;
  assign \new_Sorter100|13637_  = \new_Sorter100|13536_  | \new_Sorter100|13537_ ;
  assign \new_Sorter100|13638_  = \new_Sorter100|13538_  & \new_Sorter100|13539_ ;
  assign \new_Sorter100|13639_  = \new_Sorter100|13538_  | \new_Sorter100|13539_ ;
  assign \new_Sorter100|13640_  = \new_Sorter100|13540_  & \new_Sorter100|13541_ ;
  assign \new_Sorter100|13641_  = \new_Sorter100|13540_  | \new_Sorter100|13541_ ;
  assign \new_Sorter100|13642_  = \new_Sorter100|13542_  & \new_Sorter100|13543_ ;
  assign \new_Sorter100|13643_  = \new_Sorter100|13542_  | \new_Sorter100|13543_ ;
  assign \new_Sorter100|13644_  = \new_Sorter100|13544_  & \new_Sorter100|13545_ ;
  assign \new_Sorter100|13645_  = \new_Sorter100|13544_  | \new_Sorter100|13545_ ;
  assign \new_Sorter100|13646_  = \new_Sorter100|13546_  & \new_Sorter100|13547_ ;
  assign \new_Sorter100|13647_  = \new_Sorter100|13546_  | \new_Sorter100|13547_ ;
  assign \new_Sorter100|13648_  = \new_Sorter100|13548_  & \new_Sorter100|13549_ ;
  assign \new_Sorter100|13649_  = \new_Sorter100|13548_  | \new_Sorter100|13549_ ;
  assign \new_Sorter100|13650_  = \new_Sorter100|13550_  & \new_Sorter100|13551_ ;
  assign \new_Sorter100|13651_  = \new_Sorter100|13550_  | \new_Sorter100|13551_ ;
  assign \new_Sorter100|13652_  = \new_Sorter100|13552_  & \new_Sorter100|13553_ ;
  assign \new_Sorter100|13653_  = \new_Sorter100|13552_  | \new_Sorter100|13553_ ;
  assign \new_Sorter100|13654_  = \new_Sorter100|13554_  & \new_Sorter100|13555_ ;
  assign \new_Sorter100|13655_  = \new_Sorter100|13554_  | \new_Sorter100|13555_ ;
  assign \new_Sorter100|13656_  = \new_Sorter100|13556_  & \new_Sorter100|13557_ ;
  assign \new_Sorter100|13657_  = \new_Sorter100|13556_  | \new_Sorter100|13557_ ;
  assign \new_Sorter100|13658_  = \new_Sorter100|13558_  & \new_Sorter100|13559_ ;
  assign \new_Sorter100|13659_  = \new_Sorter100|13558_  | \new_Sorter100|13559_ ;
  assign \new_Sorter100|13660_  = \new_Sorter100|13560_  & \new_Sorter100|13561_ ;
  assign \new_Sorter100|13661_  = \new_Sorter100|13560_  | \new_Sorter100|13561_ ;
  assign \new_Sorter100|13662_  = \new_Sorter100|13562_  & \new_Sorter100|13563_ ;
  assign \new_Sorter100|13663_  = \new_Sorter100|13562_  | \new_Sorter100|13563_ ;
  assign \new_Sorter100|13664_  = \new_Sorter100|13564_  & \new_Sorter100|13565_ ;
  assign \new_Sorter100|13665_  = \new_Sorter100|13564_  | \new_Sorter100|13565_ ;
  assign \new_Sorter100|13666_  = \new_Sorter100|13566_  & \new_Sorter100|13567_ ;
  assign \new_Sorter100|13667_  = \new_Sorter100|13566_  | \new_Sorter100|13567_ ;
  assign \new_Sorter100|13668_  = \new_Sorter100|13568_  & \new_Sorter100|13569_ ;
  assign \new_Sorter100|13669_  = \new_Sorter100|13568_  | \new_Sorter100|13569_ ;
  assign \new_Sorter100|13670_  = \new_Sorter100|13570_  & \new_Sorter100|13571_ ;
  assign \new_Sorter100|13671_  = \new_Sorter100|13570_  | \new_Sorter100|13571_ ;
  assign \new_Sorter100|13672_  = \new_Sorter100|13572_  & \new_Sorter100|13573_ ;
  assign \new_Sorter100|13673_  = \new_Sorter100|13572_  | \new_Sorter100|13573_ ;
  assign \new_Sorter100|13674_  = \new_Sorter100|13574_  & \new_Sorter100|13575_ ;
  assign \new_Sorter100|13675_  = \new_Sorter100|13574_  | \new_Sorter100|13575_ ;
  assign \new_Sorter100|13676_  = \new_Sorter100|13576_  & \new_Sorter100|13577_ ;
  assign \new_Sorter100|13677_  = \new_Sorter100|13576_  | \new_Sorter100|13577_ ;
  assign \new_Sorter100|13678_  = \new_Sorter100|13578_  & \new_Sorter100|13579_ ;
  assign \new_Sorter100|13679_  = \new_Sorter100|13578_  | \new_Sorter100|13579_ ;
  assign \new_Sorter100|13680_  = \new_Sorter100|13580_  & \new_Sorter100|13581_ ;
  assign \new_Sorter100|13681_  = \new_Sorter100|13580_  | \new_Sorter100|13581_ ;
  assign \new_Sorter100|13682_  = \new_Sorter100|13582_  & \new_Sorter100|13583_ ;
  assign \new_Sorter100|13683_  = \new_Sorter100|13582_  | \new_Sorter100|13583_ ;
  assign \new_Sorter100|13684_  = \new_Sorter100|13584_  & \new_Sorter100|13585_ ;
  assign \new_Sorter100|13685_  = \new_Sorter100|13584_  | \new_Sorter100|13585_ ;
  assign \new_Sorter100|13686_  = \new_Sorter100|13586_  & \new_Sorter100|13587_ ;
  assign \new_Sorter100|13687_  = \new_Sorter100|13586_  | \new_Sorter100|13587_ ;
  assign \new_Sorter100|13688_  = \new_Sorter100|13588_  & \new_Sorter100|13589_ ;
  assign \new_Sorter100|13689_  = \new_Sorter100|13588_  | \new_Sorter100|13589_ ;
  assign \new_Sorter100|13690_  = \new_Sorter100|13590_  & \new_Sorter100|13591_ ;
  assign \new_Sorter100|13691_  = \new_Sorter100|13590_  | \new_Sorter100|13591_ ;
  assign \new_Sorter100|13692_  = \new_Sorter100|13592_  & \new_Sorter100|13593_ ;
  assign \new_Sorter100|13693_  = \new_Sorter100|13592_  | \new_Sorter100|13593_ ;
  assign \new_Sorter100|13694_  = \new_Sorter100|13594_  & \new_Sorter100|13595_ ;
  assign \new_Sorter100|13695_  = \new_Sorter100|13594_  | \new_Sorter100|13595_ ;
  assign \new_Sorter100|13696_  = \new_Sorter100|13596_  & \new_Sorter100|13597_ ;
  assign \new_Sorter100|13697_  = \new_Sorter100|13596_  | \new_Sorter100|13597_ ;
  assign \new_Sorter100|13698_  = \new_Sorter100|13598_  & \new_Sorter100|13599_ ;
  assign \new_Sorter100|13699_  = \new_Sorter100|13598_  | \new_Sorter100|13599_ ;
  assign \new_Sorter100|13700_  = \new_Sorter100|13600_ ;
  assign \new_Sorter100|13799_  = \new_Sorter100|13699_ ;
  assign \new_Sorter100|13701_  = \new_Sorter100|13601_  & \new_Sorter100|13602_ ;
  assign \new_Sorter100|13702_  = \new_Sorter100|13601_  | \new_Sorter100|13602_ ;
  assign \new_Sorter100|13703_  = \new_Sorter100|13603_  & \new_Sorter100|13604_ ;
  assign \new_Sorter100|13704_  = \new_Sorter100|13603_  | \new_Sorter100|13604_ ;
  assign \new_Sorter100|13705_  = \new_Sorter100|13605_  & \new_Sorter100|13606_ ;
  assign \new_Sorter100|13706_  = \new_Sorter100|13605_  | \new_Sorter100|13606_ ;
  assign \new_Sorter100|13707_  = \new_Sorter100|13607_  & \new_Sorter100|13608_ ;
  assign \new_Sorter100|13708_  = \new_Sorter100|13607_  | \new_Sorter100|13608_ ;
  assign \new_Sorter100|13709_  = \new_Sorter100|13609_  & \new_Sorter100|13610_ ;
  assign \new_Sorter100|13710_  = \new_Sorter100|13609_  | \new_Sorter100|13610_ ;
  assign \new_Sorter100|13711_  = \new_Sorter100|13611_  & \new_Sorter100|13612_ ;
  assign \new_Sorter100|13712_  = \new_Sorter100|13611_  | \new_Sorter100|13612_ ;
  assign \new_Sorter100|13713_  = \new_Sorter100|13613_  & \new_Sorter100|13614_ ;
  assign \new_Sorter100|13714_  = \new_Sorter100|13613_  | \new_Sorter100|13614_ ;
  assign \new_Sorter100|13715_  = \new_Sorter100|13615_  & \new_Sorter100|13616_ ;
  assign \new_Sorter100|13716_  = \new_Sorter100|13615_  | \new_Sorter100|13616_ ;
  assign \new_Sorter100|13717_  = \new_Sorter100|13617_  & \new_Sorter100|13618_ ;
  assign \new_Sorter100|13718_  = \new_Sorter100|13617_  | \new_Sorter100|13618_ ;
  assign \new_Sorter100|13719_  = \new_Sorter100|13619_  & \new_Sorter100|13620_ ;
  assign \new_Sorter100|13720_  = \new_Sorter100|13619_  | \new_Sorter100|13620_ ;
  assign \new_Sorter100|13721_  = \new_Sorter100|13621_  & \new_Sorter100|13622_ ;
  assign \new_Sorter100|13722_  = \new_Sorter100|13621_  | \new_Sorter100|13622_ ;
  assign \new_Sorter100|13723_  = \new_Sorter100|13623_  & \new_Sorter100|13624_ ;
  assign \new_Sorter100|13724_  = \new_Sorter100|13623_  | \new_Sorter100|13624_ ;
  assign \new_Sorter100|13725_  = \new_Sorter100|13625_  & \new_Sorter100|13626_ ;
  assign \new_Sorter100|13726_  = \new_Sorter100|13625_  | \new_Sorter100|13626_ ;
  assign \new_Sorter100|13727_  = \new_Sorter100|13627_  & \new_Sorter100|13628_ ;
  assign \new_Sorter100|13728_  = \new_Sorter100|13627_  | \new_Sorter100|13628_ ;
  assign \new_Sorter100|13729_  = \new_Sorter100|13629_  & \new_Sorter100|13630_ ;
  assign \new_Sorter100|13730_  = \new_Sorter100|13629_  | \new_Sorter100|13630_ ;
  assign \new_Sorter100|13731_  = \new_Sorter100|13631_  & \new_Sorter100|13632_ ;
  assign \new_Sorter100|13732_  = \new_Sorter100|13631_  | \new_Sorter100|13632_ ;
  assign \new_Sorter100|13733_  = \new_Sorter100|13633_  & \new_Sorter100|13634_ ;
  assign \new_Sorter100|13734_  = \new_Sorter100|13633_  | \new_Sorter100|13634_ ;
  assign \new_Sorter100|13735_  = \new_Sorter100|13635_  & \new_Sorter100|13636_ ;
  assign \new_Sorter100|13736_  = \new_Sorter100|13635_  | \new_Sorter100|13636_ ;
  assign \new_Sorter100|13737_  = \new_Sorter100|13637_  & \new_Sorter100|13638_ ;
  assign \new_Sorter100|13738_  = \new_Sorter100|13637_  | \new_Sorter100|13638_ ;
  assign \new_Sorter100|13739_  = \new_Sorter100|13639_  & \new_Sorter100|13640_ ;
  assign \new_Sorter100|13740_  = \new_Sorter100|13639_  | \new_Sorter100|13640_ ;
  assign \new_Sorter100|13741_  = \new_Sorter100|13641_  & \new_Sorter100|13642_ ;
  assign \new_Sorter100|13742_  = \new_Sorter100|13641_  | \new_Sorter100|13642_ ;
  assign \new_Sorter100|13743_  = \new_Sorter100|13643_  & \new_Sorter100|13644_ ;
  assign \new_Sorter100|13744_  = \new_Sorter100|13643_  | \new_Sorter100|13644_ ;
  assign \new_Sorter100|13745_  = \new_Sorter100|13645_  & \new_Sorter100|13646_ ;
  assign \new_Sorter100|13746_  = \new_Sorter100|13645_  | \new_Sorter100|13646_ ;
  assign \new_Sorter100|13747_  = \new_Sorter100|13647_  & \new_Sorter100|13648_ ;
  assign \new_Sorter100|13748_  = \new_Sorter100|13647_  | \new_Sorter100|13648_ ;
  assign \new_Sorter100|13749_  = \new_Sorter100|13649_  & \new_Sorter100|13650_ ;
  assign \new_Sorter100|13750_  = \new_Sorter100|13649_  | \new_Sorter100|13650_ ;
  assign \new_Sorter100|13751_  = \new_Sorter100|13651_  & \new_Sorter100|13652_ ;
  assign \new_Sorter100|13752_  = \new_Sorter100|13651_  | \new_Sorter100|13652_ ;
  assign \new_Sorter100|13753_  = \new_Sorter100|13653_  & \new_Sorter100|13654_ ;
  assign \new_Sorter100|13754_  = \new_Sorter100|13653_  | \new_Sorter100|13654_ ;
  assign \new_Sorter100|13755_  = \new_Sorter100|13655_  & \new_Sorter100|13656_ ;
  assign \new_Sorter100|13756_  = \new_Sorter100|13655_  | \new_Sorter100|13656_ ;
  assign \new_Sorter100|13757_  = \new_Sorter100|13657_  & \new_Sorter100|13658_ ;
  assign \new_Sorter100|13758_  = \new_Sorter100|13657_  | \new_Sorter100|13658_ ;
  assign \new_Sorter100|13759_  = \new_Sorter100|13659_  & \new_Sorter100|13660_ ;
  assign \new_Sorter100|13760_  = \new_Sorter100|13659_  | \new_Sorter100|13660_ ;
  assign \new_Sorter100|13761_  = \new_Sorter100|13661_  & \new_Sorter100|13662_ ;
  assign \new_Sorter100|13762_  = \new_Sorter100|13661_  | \new_Sorter100|13662_ ;
  assign \new_Sorter100|13763_  = \new_Sorter100|13663_  & \new_Sorter100|13664_ ;
  assign \new_Sorter100|13764_  = \new_Sorter100|13663_  | \new_Sorter100|13664_ ;
  assign \new_Sorter100|13765_  = \new_Sorter100|13665_  & \new_Sorter100|13666_ ;
  assign \new_Sorter100|13766_  = \new_Sorter100|13665_  | \new_Sorter100|13666_ ;
  assign \new_Sorter100|13767_  = \new_Sorter100|13667_  & \new_Sorter100|13668_ ;
  assign \new_Sorter100|13768_  = \new_Sorter100|13667_  | \new_Sorter100|13668_ ;
  assign \new_Sorter100|13769_  = \new_Sorter100|13669_  & \new_Sorter100|13670_ ;
  assign \new_Sorter100|13770_  = \new_Sorter100|13669_  | \new_Sorter100|13670_ ;
  assign \new_Sorter100|13771_  = \new_Sorter100|13671_  & \new_Sorter100|13672_ ;
  assign \new_Sorter100|13772_  = \new_Sorter100|13671_  | \new_Sorter100|13672_ ;
  assign \new_Sorter100|13773_  = \new_Sorter100|13673_  & \new_Sorter100|13674_ ;
  assign \new_Sorter100|13774_  = \new_Sorter100|13673_  | \new_Sorter100|13674_ ;
  assign \new_Sorter100|13775_  = \new_Sorter100|13675_  & \new_Sorter100|13676_ ;
  assign \new_Sorter100|13776_  = \new_Sorter100|13675_  | \new_Sorter100|13676_ ;
  assign \new_Sorter100|13777_  = \new_Sorter100|13677_  & \new_Sorter100|13678_ ;
  assign \new_Sorter100|13778_  = \new_Sorter100|13677_  | \new_Sorter100|13678_ ;
  assign \new_Sorter100|13779_  = \new_Sorter100|13679_  & \new_Sorter100|13680_ ;
  assign \new_Sorter100|13780_  = \new_Sorter100|13679_  | \new_Sorter100|13680_ ;
  assign \new_Sorter100|13781_  = \new_Sorter100|13681_  & \new_Sorter100|13682_ ;
  assign \new_Sorter100|13782_  = \new_Sorter100|13681_  | \new_Sorter100|13682_ ;
  assign \new_Sorter100|13783_  = \new_Sorter100|13683_  & \new_Sorter100|13684_ ;
  assign \new_Sorter100|13784_  = \new_Sorter100|13683_  | \new_Sorter100|13684_ ;
  assign \new_Sorter100|13785_  = \new_Sorter100|13685_  & \new_Sorter100|13686_ ;
  assign \new_Sorter100|13786_  = \new_Sorter100|13685_  | \new_Sorter100|13686_ ;
  assign \new_Sorter100|13787_  = \new_Sorter100|13687_  & \new_Sorter100|13688_ ;
  assign \new_Sorter100|13788_  = \new_Sorter100|13687_  | \new_Sorter100|13688_ ;
  assign \new_Sorter100|13789_  = \new_Sorter100|13689_  & \new_Sorter100|13690_ ;
  assign \new_Sorter100|13790_  = \new_Sorter100|13689_  | \new_Sorter100|13690_ ;
  assign \new_Sorter100|13791_  = \new_Sorter100|13691_  & \new_Sorter100|13692_ ;
  assign \new_Sorter100|13792_  = \new_Sorter100|13691_  | \new_Sorter100|13692_ ;
  assign \new_Sorter100|13793_  = \new_Sorter100|13693_  & \new_Sorter100|13694_ ;
  assign \new_Sorter100|13794_  = \new_Sorter100|13693_  | \new_Sorter100|13694_ ;
  assign \new_Sorter100|13795_  = \new_Sorter100|13695_  & \new_Sorter100|13696_ ;
  assign \new_Sorter100|13796_  = \new_Sorter100|13695_  | \new_Sorter100|13696_ ;
  assign \new_Sorter100|13797_  = \new_Sorter100|13697_  & \new_Sorter100|13698_ ;
  assign \new_Sorter100|13798_  = \new_Sorter100|13697_  | \new_Sorter100|13698_ ;
  assign \new_Sorter100|13800_  = \new_Sorter100|13700_  & \new_Sorter100|13701_ ;
  assign \new_Sorter100|13801_  = \new_Sorter100|13700_  | \new_Sorter100|13701_ ;
  assign \new_Sorter100|13802_  = \new_Sorter100|13702_  & \new_Sorter100|13703_ ;
  assign \new_Sorter100|13803_  = \new_Sorter100|13702_  | \new_Sorter100|13703_ ;
  assign \new_Sorter100|13804_  = \new_Sorter100|13704_  & \new_Sorter100|13705_ ;
  assign \new_Sorter100|13805_  = \new_Sorter100|13704_  | \new_Sorter100|13705_ ;
  assign \new_Sorter100|13806_  = \new_Sorter100|13706_  & \new_Sorter100|13707_ ;
  assign \new_Sorter100|13807_  = \new_Sorter100|13706_  | \new_Sorter100|13707_ ;
  assign \new_Sorter100|13808_  = \new_Sorter100|13708_  & \new_Sorter100|13709_ ;
  assign \new_Sorter100|13809_  = \new_Sorter100|13708_  | \new_Sorter100|13709_ ;
  assign \new_Sorter100|13810_  = \new_Sorter100|13710_  & \new_Sorter100|13711_ ;
  assign \new_Sorter100|13811_  = \new_Sorter100|13710_  | \new_Sorter100|13711_ ;
  assign \new_Sorter100|13812_  = \new_Sorter100|13712_  & \new_Sorter100|13713_ ;
  assign \new_Sorter100|13813_  = \new_Sorter100|13712_  | \new_Sorter100|13713_ ;
  assign \new_Sorter100|13814_  = \new_Sorter100|13714_  & \new_Sorter100|13715_ ;
  assign \new_Sorter100|13815_  = \new_Sorter100|13714_  | \new_Sorter100|13715_ ;
  assign \new_Sorter100|13816_  = \new_Sorter100|13716_  & \new_Sorter100|13717_ ;
  assign \new_Sorter100|13817_  = \new_Sorter100|13716_  | \new_Sorter100|13717_ ;
  assign \new_Sorter100|13818_  = \new_Sorter100|13718_  & \new_Sorter100|13719_ ;
  assign \new_Sorter100|13819_  = \new_Sorter100|13718_  | \new_Sorter100|13719_ ;
  assign \new_Sorter100|13820_  = \new_Sorter100|13720_  & \new_Sorter100|13721_ ;
  assign \new_Sorter100|13821_  = \new_Sorter100|13720_  | \new_Sorter100|13721_ ;
  assign \new_Sorter100|13822_  = \new_Sorter100|13722_  & \new_Sorter100|13723_ ;
  assign \new_Sorter100|13823_  = \new_Sorter100|13722_  | \new_Sorter100|13723_ ;
  assign \new_Sorter100|13824_  = \new_Sorter100|13724_  & \new_Sorter100|13725_ ;
  assign \new_Sorter100|13825_  = \new_Sorter100|13724_  | \new_Sorter100|13725_ ;
  assign \new_Sorter100|13826_  = \new_Sorter100|13726_  & \new_Sorter100|13727_ ;
  assign \new_Sorter100|13827_  = \new_Sorter100|13726_  | \new_Sorter100|13727_ ;
  assign \new_Sorter100|13828_  = \new_Sorter100|13728_  & \new_Sorter100|13729_ ;
  assign \new_Sorter100|13829_  = \new_Sorter100|13728_  | \new_Sorter100|13729_ ;
  assign \new_Sorter100|13830_  = \new_Sorter100|13730_  & \new_Sorter100|13731_ ;
  assign \new_Sorter100|13831_  = \new_Sorter100|13730_  | \new_Sorter100|13731_ ;
  assign \new_Sorter100|13832_  = \new_Sorter100|13732_  & \new_Sorter100|13733_ ;
  assign \new_Sorter100|13833_  = \new_Sorter100|13732_  | \new_Sorter100|13733_ ;
  assign \new_Sorter100|13834_  = \new_Sorter100|13734_  & \new_Sorter100|13735_ ;
  assign \new_Sorter100|13835_  = \new_Sorter100|13734_  | \new_Sorter100|13735_ ;
  assign \new_Sorter100|13836_  = \new_Sorter100|13736_  & \new_Sorter100|13737_ ;
  assign \new_Sorter100|13837_  = \new_Sorter100|13736_  | \new_Sorter100|13737_ ;
  assign \new_Sorter100|13838_  = \new_Sorter100|13738_  & \new_Sorter100|13739_ ;
  assign \new_Sorter100|13839_  = \new_Sorter100|13738_  | \new_Sorter100|13739_ ;
  assign \new_Sorter100|13840_  = \new_Sorter100|13740_  & \new_Sorter100|13741_ ;
  assign \new_Sorter100|13841_  = \new_Sorter100|13740_  | \new_Sorter100|13741_ ;
  assign \new_Sorter100|13842_  = \new_Sorter100|13742_  & \new_Sorter100|13743_ ;
  assign \new_Sorter100|13843_  = \new_Sorter100|13742_  | \new_Sorter100|13743_ ;
  assign \new_Sorter100|13844_  = \new_Sorter100|13744_  & \new_Sorter100|13745_ ;
  assign \new_Sorter100|13845_  = \new_Sorter100|13744_  | \new_Sorter100|13745_ ;
  assign \new_Sorter100|13846_  = \new_Sorter100|13746_  & \new_Sorter100|13747_ ;
  assign \new_Sorter100|13847_  = \new_Sorter100|13746_  | \new_Sorter100|13747_ ;
  assign \new_Sorter100|13848_  = \new_Sorter100|13748_  & \new_Sorter100|13749_ ;
  assign \new_Sorter100|13849_  = \new_Sorter100|13748_  | \new_Sorter100|13749_ ;
  assign \new_Sorter100|13850_  = \new_Sorter100|13750_  & \new_Sorter100|13751_ ;
  assign \new_Sorter100|13851_  = \new_Sorter100|13750_  | \new_Sorter100|13751_ ;
  assign \new_Sorter100|13852_  = \new_Sorter100|13752_  & \new_Sorter100|13753_ ;
  assign \new_Sorter100|13853_  = \new_Sorter100|13752_  | \new_Sorter100|13753_ ;
  assign \new_Sorter100|13854_  = \new_Sorter100|13754_  & \new_Sorter100|13755_ ;
  assign \new_Sorter100|13855_  = \new_Sorter100|13754_  | \new_Sorter100|13755_ ;
  assign \new_Sorter100|13856_  = \new_Sorter100|13756_  & \new_Sorter100|13757_ ;
  assign \new_Sorter100|13857_  = \new_Sorter100|13756_  | \new_Sorter100|13757_ ;
  assign \new_Sorter100|13858_  = \new_Sorter100|13758_  & \new_Sorter100|13759_ ;
  assign \new_Sorter100|13859_  = \new_Sorter100|13758_  | \new_Sorter100|13759_ ;
  assign \new_Sorter100|13860_  = \new_Sorter100|13760_  & \new_Sorter100|13761_ ;
  assign \new_Sorter100|13861_  = \new_Sorter100|13760_  | \new_Sorter100|13761_ ;
  assign \new_Sorter100|13862_  = \new_Sorter100|13762_  & \new_Sorter100|13763_ ;
  assign \new_Sorter100|13863_  = \new_Sorter100|13762_  | \new_Sorter100|13763_ ;
  assign \new_Sorter100|13864_  = \new_Sorter100|13764_  & \new_Sorter100|13765_ ;
  assign \new_Sorter100|13865_  = \new_Sorter100|13764_  | \new_Sorter100|13765_ ;
  assign \new_Sorter100|13866_  = \new_Sorter100|13766_  & \new_Sorter100|13767_ ;
  assign \new_Sorter100|13867_  = \new_Sorter100|13766_  | \new_Sorter100|13767_ ;
  assign \new_Sorter100|13868_  = \new_Sorter100|13768_  & \new_Sorter100|13769_ ;
  assign \new_Sorter100|13869_  = \new_Sorter100|13768_  | \new_Sorter100|13769_ ;
  assign \new_Sorter100|13870_  = \new_Sorter100|13770_  & \new_Sorter100|13771_ ;
  assign \new_Sorter100|13871_  = \new_Sorter100|13770_  | \new_Sorter100|13771_ ;
  assign \new_Sorter100|13872_  = \new_Sorter100|13772_  & \new_Sorter100|13773_ ;
  assign \new_Sorter100|13873_  = \new_Sorter100|13772_  | \new_Sorter100|13773_ ;
  assign \new_Sorter100|13874_  = \new_Sorter100|13774_  & \new_Sorter100|13775_ ;
  assign \new_Sorter100|13875_  = \new_Sorter100|13774_  | \new_Sorter100|13775_ ;
  assign \new_Sorter100|13876_  = \new_Sorter100|13776_  & \new_Sorter100|13777_ ;
  assign \new_Sorter100|13877_  = \new_Sorter100|13776_  | \new_Sorter100|13777_ ;
  assign \new_Sorter100|13878_  = \new_Sorter100|13778_  & \new_Sorter100|13779_ ;
  assign \new_Sorter100|13879_  = \new_Sorter100|13778_  | \new_Sorter100|13779_ ;
  assign \new_Sorter100|13880_  = \new_Sorter100|13780_  & \new_Sorter100|13781_ ;
  assign \new_Sorter100|13881_  = \new_Sorter100|13780_  | \new_Sorter100|13781_ ;
  assign \new_Sorter100|13882_  = \new_Sorter100|13782_  & \new_Sorter100|13783_ ;
  assign \new_Sorter100|13883_  = \new_Sorter100|13782_  | \new_Sorter100|13783_ ;
  assign \new_Sorter100|13884_  = \new_Sorter100|13784_  & \new_Sorter100|13785_ ;
  assign \new_Sorter100|13885_  = \new_Sorter100|13784_  | \new_Sorter100|13785_ ;
  assign \new_Sorter100|13886_  = \new_Sorter100|13786_  & \new_Sorter100|13787_ ;
  assign \new_Sorter100|13887_  = \new_Sorter100|13786_  | \new_Sorter100|13787_ ;
  assign \new_Sorter100|13888_  = \new_Sorter100|13788_  & \new_Sorter100|13789_ ;
  assign \new_Sorter100|13889_  = \new_Sorter100|13788_  | \new_Sorter100|13789_ ;
  assign \new_Sorter100|13890_  = \new_Sorter100|13790_  & \new_Sorter100|13791_ ;
  assign \new_Sorter100|13891_  = \new_Sorter100|13790_  | \new_Sorter100|13791_ ;
  assign \new_Sorter100|13892_  = \new_Sorter100|13792_  & \new_Sorter100|13793_ ;
  assign \new_Sorter100|13893_  = \new_Sorter100|13792_  | \new_Sorter100|13793_ ;
  assign \new_Sorter100|13894_  = \new_Sorter100|13794_  & \new_Sorter100|13795_ ;
  assign \new_Sorter100|13895_  = \new_Sorter100|13794_  | \new_Sorter100|13795_ ;
  assign \new_Sorter100|13896_  = \new_Sorter100|13796_  & \new_Sorter100|13797_ ;
  assign \new_Sorter100|13897_  = \new_Sorter100|13796_  | \new_Sorter100|13797_ ;
  assign \new_Sorter100|13898_  = \new_Sorter100|13798_  & \new_Sorter100|13799_ ;
  assign \new_Sorter100|13899_  = \new_Sorter100|13798_  | \new_Sorter100|13799_ ;
  assign \new_Sorter100|13900_  = \new_Sorter100|13800_ ;
  assign \new_Sorter100|13999_  = \new_Sorter100|13899_ ;
  assign \new_Sorter100|13901_  = \new_Sorter100|13801_  & \new_Sorter100|13802_ ;
  assign \new_Sorter100|13902_  = \new_Sorter100|13801_  | \new_Sorter100|13802_ ;
  assign \new_Sorter100|13903_  = \new_Sorter100|13803_  & \new_Sorter100|13804_ ;
  assign \new_Sorter100|13904_  = \new_Sorter100|13803_  | \new_Sorter100|13804_ ;
  assign \new_Sorter100|13905_  = \new_Sorter100|13805_  & \new_Sorter100|13806_ ;
  assign \new_Sorter100|13906_  = \new_Sorter100|13805_  | \new_Sorter100|13806_ ;
  assign \new_Sorter100|13907_  = \new_Sorter100|13807_  & \new_Sorter100|13808_ ;
  assign \new_Sorter100|13908_  = \new_Sorter100|13807_  | \new_Sorter100|13808_ ;
  assign \new_Sorter100|13909_  = \new_Sorter100|13809_  & \new_Sorter100|13810_ ;
  assign \new_Sorter100|13910_  = \new_Sorter100|13809_  | \new_Sorter100|13810_ ;
  assign \new_Sorter100|13911_  = \new_Sorter100|13811_  & \new_Sorter100|13812_ ;
  assign \new_Sorter100|13912_  = \new_Sorter100|13811_  | \new_Sorter100|13812_ ;
  assign \new_Sorter100|13913_  = \new_Sorter100|13813_  & \new_Sorter100|13814_ ;
  assign \new_Sorter100|13914_  = \new_Sorter100|13813_  | \new_Sorter100|13814_ ;
  assign \new_Sorter100|13915_  = \new_Sorter100|13815_  & \new_Sorter100|13816_ ;
  assign \new_Sorter100|13916_  = \new_Sorter100|13815_  | \new_Sorter100|13816_ ;
  assign \new_Sorter100|13917_  = \new_Sorter100|13817_  & \new_Sorter100|13818_ ;
  assign \new_Sorter100|13918_  = \new_Sorter100|13817_  | \new_Sorter100|13818_ ;
  assign \new_Sorter100|13919_  = \new_Sorter100|13819_  & \new_Sorter100|13820_ ;
  assign \new_Sorter100|13920_  = \new_Sorter100|13819_  | \new_Sorter100|13820_ ;
  assign \new_Sorter100|13921_  = \new_Sorter100|13821_  & \new_Sorter100|13822_ ;
  assign \new_Sorter100|13922_  = \new_Sorter100|13821_  | \new_Sorter100|13822_ ;
  assign \new_Sorter100|13923_  = \new_Sorter100|13823_  & \new_Sorter100|13824_ ;
  assign \new_Sorter100|13924_  = \new_Sorter100|13823_  | \new_Sorter100|13824_ ;
  assign \new_Sorter100|13925_  = \new_Sorter100|13825_  & \new_Sorter100|13826_ ;
  assign \new_Sorter100|13926_  = \new_Sorter100|13825_  | \new_Sorter100|13826_ ;
  assign \new_Sorter100|13927_  = \new_Sorter100|13827_  & \new_Sorter100|13828_ ;
  assign \new_Sorter100|13928_  = \new_Sorter100|13827_  | \new_Sorter100|13828_ ;
  assign \new_Sorter100|13929_  = \new_Sorter100|13829_  & \new_Sorter100|13830_ ;
  assign \new_Sorter100|13930_  = \new_Sorter100|13829_  | \new_Sorter100|13830_ ;
  assign \new_Sorter100|13931_  = \new_Sorter100|13831_  & \new_Sorter100|13832_ ;
  assign \new_Sorter100|13932_  = \new_Sorter100|13831_  | \new_Sorter100|13832_ ;
  assign \new_Sorter100|13933_  = \new_Sorter100|13833_  & \new_Sorter100|13834_ ;
  assign \new_Sorter100|13934_  = \new_Sorter100|13833_  | \new_Sorter100|13834_ ;
  assign \new_Sorter100|13935_  = \new_Sorter100|13835_  & \new_Sorter100|13836_ ;
  assign \new_Sorter100|13936_  = \new_Sorter100|13835_  | \new_Sorter100|13836_ ;
  assign \new_Sorter100|13937_  = \new_Sorter100|13837_  & \new_Sorter100|13838_ ;
  assign \new_Sorter100|13938_  = \new_Sorter100|13837_  | \new_Sorter100|13838_ ;
  assign \new_Sorter100|13939_  = \new_Sorter100|13839_  & \new_Sorter100|13840_ ;
  assign \new_Sorter100|13940_  = \new_Sorter100|13839_  | \new_Sorter100|13840_ ;
  assign \new_Sorter100|13941_  = \new_Sorter100|13841_  & \new_Sorter100|13842_ ;
  assign \new_Sorter100|13942_  = \new_Sorter100|13841_  | \new_Sorter100|13842_ ;
  assign \new_Sorter100|13943_  = \new_Sorter100|13843_  & \new_Sorter100|13844_ ;
  assign \new_Sorter100|13944_  = \new_Sorter100|13843_  | \new_Sorter100|13844_ ;
  assign \new_Sorter100|13945_  = \new_Sorter100|13845_  & \new_Sorter100|13846_ ;
  assign \new_Sorter100|13946_  = \new_Sorter100|13845_  | \new_Sorter100|13846_ ;
  assign \new_Sorter100|13947_  = \new_Sorter100|13847_  & \new_Sorter100|13848_ ;
  assign \new_Sorter100|13948_  = \new_Sorter100|13847_  | \new_Sorter100|13848_ ;
  assign \new_Sorter100|13949_  = \new_Sorter100|13849_  & \new_Sorter100|13850_ ;
  assign \new_Sorter100|13950_  = \new_Sorter100|13849_  | \new_Sorter100|13850_ ;
  assign \new_Sorter100|13951_  = \new_Sorter100|13851_  & \new_Sorter100|13852_ ;
  assign \new_Sorter100|13952_  = \new_Sorter100|13851_  | \new_Sorter100|13852_ ;
  assign \new_Sorter100|13953_  = \new_Sorter100|13853_  & \new_Sorter100|13854_ ;
  assign \new_Sorter100|13954_  = \new_Sorter100|13853_  | \new_Sorter100|13854_ ;
  assign \new_Sorter100|13955_  = \new_Sorter100|13855_  & \new_Sorter100|13856_ ;
  assign \new_Sorter100|13956_  = \new_Sorter100|13855_  | \new_Sorter100|13856_ ;
  assign \new_Sorter100|13957_  = \new_Sorter100|13857_  & \new_Sorter100|13858_ ;
  assign \new_Sorter100|13958_  = \new_Sorter100|13857_  | \new_Sorter100|13858_ ;
  assign \new_Sorter100|13959_  = \new_Sorter100|13859_  & \new_Sorter100|13860_ ;
  assign \new_Sorter100|13960_  = \new_Sorter100|13859_  | \new_Sorter100|13860_ ;
  assign \new_Sorter100|13961_  = \new_Sorter100|13861_  & \new_Sorter100|13862_ ;
  assign \new_Sorter100|13962_  = \new_Sorter100|13861_  | \new_Sorter100|13862_ ;
  assign \new_Sorter100|13963_  = \new_Sorter100|13863_  & \new_Sorter100|13864_ ;
  assign \new_Sorter100|13964_  = \new_Sorter100|13863_  | \new_Sorter100|13864_ ;
  assign \new_Sorter100|13965_  = \new_Sorter100|13865_  & \new_Sorter100|13866_ ;
  assign \new_Sorter100|13966_  = \new_Sorter100|13865_  | \new_Sorter100|13866_ ;
  assign \new_Sorter100|13967_  = \new_Sorter100|13867_  & \new_Sorter100|13868_ ;
  assign \new_Sorter100|13968_  = \new_Sorter100|13867_  | \new_Sorter100|13868_ ;
  assign \new_Sorter100|13969_  = \new_Sorter100|13869_  & \new_Sorter100|13870_ ;
  assign \new_Sorter100|13970_  = \new_Sorter100|13869_  | \new_Sorter100|13870_ ;
  assign \new_Sorter100|13971_  = \new_Sorter100|13871_  & \new_Sorter100|13872_ ;
  assign \new_Sorter100|13972_  = \new_Sorter100|13871_  | \new_Sorter100|13872_ ;
  assign \new_Sorter100|13973_  = \new_Sorter100|13873_  & \new_Sorter100|13874_ ;
  assign \new_Sorter100|13974_  = \new_Sorter100|13873_  | \new_Sorter100|13874_ ;
  assign \new_Sorter100|13975_  = \new_Sorter100|13875_  & \new_Sorter100|13876_ ;
  assign \new_Sorter100|13976_  = \new_Sorter100|13875_  | \new_Sorter100|13876_ ;
  assign \new_Sorter100|13977_  = \new_Sorter100|13877_  & \new_Sorter100|13878_ ;
  assign \new_Sorter100|13978_  = \new_Sorter100|13877_  | \new_Sorter100|13878_ ;
  assign \new_Sorter100|13979_  = \new_Sorter100|13879_  & \new_Sorter100|13880_ ;
  assign \new_Sorter100|13980_  = \new_Sorter100|13879_  | \new_Sorter100|13880_ ;
  assign \new_Sorter100|13981_  = \new_Sorter100|13881_  & \new_Sorter100|13882_ ;
  assign \new_Sorter100|13982_  = \new_Sorter100|13881_  | \new_Sorter100|13882_ ;
  assign \new_Sorter100|13983_  = \new_Sorter100|13883_  & \new_Sorter100|13884_ ;
  assign \new_Sorter100|13984_  = \new_Sorter100|13883_  | \new_Sorter100|13884_ ;
  assign \new_Sorter100|13985_  = \new_Sorter100|13885_  & \new_Sorter100|13886_ ;
  assign \new_Sorter100|13986_  = \new_Sorter100|13885_  | \new_Sorter100|13886_ ;
  assign \new_Sorter100|13987_  = \new_Sorter100|13887_  & \new_Sorter100|13888_ ;
  assign \new_Sorter100|13988_  = \new_Sorter100|13887_  | \new_Sorter100|13888_ ;
  assign \new_Sorter100|13989_  = \new_Sorter100|13889_  & \new_Sorter100|13890_ ;
  assign \new_Sorter100|13990_  = \new_Sorter100|13889_  | \new_Sorter100|13890_ ;
  assign \new_Sorter100|13991_  = \new_Sorter100|13891_  & \new_Sorter100|13892_ ;
  assign \new_Sorter100|13992_  = \new_Sorter100|13891_  | \new_Sorter100|13892_ ;
  assign \new_Sorter100|13993_  = \new_Sorter100|13893_  & \new_Sorter100|13894_ ;
  assign \new_Sorter100|13994_  = \new_Sorter100|13893_  | \new_Sorter100|13894_ ;
  assign \new_Sorter100|13995_  = \new_Sorter100|13895_  & \new_Sorter100|13896_ ;
  assign \new_Sorter100|13996_  = \new_Sorter100|13895_  | \new_Sorter100|13896_ ;
  assign \new_Sorter100|13997_  = \new_Sorter100|13897_  & \new_Sorter100|13898_ ;
  assign \new_Sorter100|13998_  = \new_Sorter100|13897_  | \new_Sorter100|13898_ ;
  assign \new_Sorter100|14000_  = \new_Sorter100|13900_  & \new_Sorter100|13901_ ;
  assign \new_Sorter100|14001_  = \new_Sorter100|13900_  | \new_Sorter100|13901_ ;
  assign \new_Sorter100|14002_  = \new_Sorter100|13902_  & \new_Sorter100|13903_ ;
  assign \new_Sorter100|14003_  = \new_Sorter100|13902_  | \new_Sorter100|13903_ ;
  assign \new_Sorter100|14004_  = \new_Sorter100|13904_  & \new_Sorter100|13905_ ;
  assign \new_Sorter100|14005_  = \new_Sorter100|13904_  | \new_Sorter100|13905_ ;
  assign \new_Sorter100|14006_  = \new_Sorter100|13906_  & \new_Sorter100|13907_ ;
  assign \new_Sorter100|14007_  = \new_Sorter100|13906_  | \new_Sorter100|13907_ ;
  assign \new_Sorter100|14008_  = \new_Sorter100|13908_  & \new_Sorter100|13909_ ;
  assign \new_Sorter100|14009_  = \new_Sorter100|13908_  | \new_Sorter100|13909_ ;
  assign \new_Sorter100|14010_  = \new_Sorter100|13910_  & \new_Sorter100|13911_ ;
  assign \new_Sorter100|14011_  = \new_Sorter100|13910_  | \new_Sorter100|13911_ ;
  assign \new_Sorter100|14012_  = \new_Sorter100|13912_  & \new_Sorter100|13913_ ;
  assign \new_Sorter100|14013_  = \new_Sorter100|13912_  | \new_Sorter100|13913_ ;
  assign \new_Sorter100|14014_  = \new_Sorter100|13914_  & \new_Sorter100|13915_ ;
  assign \new_Sorter100|14015_  = \new_Sorter100|13914_  | \new_Sorter100|13915_ ;
  assign \new_Sorter100|14016_  = \new_Sorter100|13916_  & \new_Sorter100|13917_ ;
  assign \new_Sorter100|14017_  = \new_Sorter100|13916_  | \new_Sorter100|13917_ ;
  assign \new_Sorter100|14018_  = \new_Sorter100|13918_  & \new_Sorter100|13919_ ;
  assign \new_Sorter100|14019_  = \new_Sorter100|13918_  | \new_Sorter100|13919_ ;
  assign \new_Sorter100|14020_  = \new_Sorter100|13920_  & \new_Sorter100|13921_ ;
  assign \new_Sorter100|14021_  = \new_Sorter100|13920_  | \new_Sorter100|13921_ ;
  assign \new_Sorter100|14022_  = \new_Sorter100|13922_  & \new_Sorter100|13923_ ;
  assign \new_Sorter100|14023_  = \new_Sorter100|13922_  | \new_Sorter100|13923_ ;
  assign \new_Sorter100|14024_  = \new_Sorter100|13924_  & \new_Sorter100|13925_ ;
  assign \new_Sorter100|14025_  = \new_Sorter100|13924_  | \new_Sorter100|13925_ ;
  assign \new_Sorter100|14026_  = \new_Sorter100|13926_  & \new_Sorter100|13927_ ;
  assign \new_Sorter100|14027_  = \new_Sorter100|13926_  | \new_Sorter100|13927_ ;
  assign \new_Sorter100|14028_  = \new_Sorter100|13928_  & \new_Sorter100|13929_ ;
  assign \new_Sorter100|14029_  = \new_Sorter100|13928_  | \new_Sorter100|13929_ ;
  assign \new_Sorter100|14030_  = \new_Sorter100|13930_  & \new_Sorter100|13931_ ;
  assign \new_Sorter100|14031_  = \new_Sorter100|13930_  | \new_Sorter100|13931_ ;
  assign \new_Sorter100|14032_  = \new_Sorter100|13932_  & \new_Sorter100|13933_ ;
  assign \new_Sorter100|14033_  = \new_Sorter100|13932_  | \new_Sorter100|13933_ ;
  assign \new_Sorter100|14034_  = \new_Sorter100|13934_  & \new_Sorter100|13935_ ;
  assign \new_Sorter100|14035_  = \new_Sorter100|13934_  | \new_Sorter100|13935_ ;
  assign \new_Sorter100|14036_  = \new_Sorter100|13936_  & \new_Sorter100|13937_ ;
  assign \new_Sorter100|14037_  = \new_Sorter100|13936_  | \new_Sorter100|13937_ ;
  assign \new_Sorter100|14038_  = \new_Sorter100|13938_  & \new_Sorter100|13939_ ;
  assign \new_Sorter100|14039_  = \new_Sorter100|13938_  | \new_Sorter100|13939_ ;
  assign \new_Sorter100|14040_  = \new_Sorter100|13940_  & \new_Sorter100|13941_ ;
  assign \new_Sorter100|14041_  = \new_Sorter100|13940_  | \new_Sorter100|13941_ ;
  assign \new_Sorter100|14042_  = \new_Sorter100|13942_  & \new_Sorter100|13943_ ;
  assign \new_Sorter100|14043_  = \new_Sorter100|13942_  | \new_Sorter100|13943_ ;
  assign \new_Sorter100|14044_  = \new_Sorter100|13944_  & \new_Sorter100|13945_ ;
  assign \new_Sorter100|14045_  = \new_Sorter100|13944_  | \new_Sorter100|13945_ ;
  assign \new_Sorter100|14046_  = \new_Sorter100|13946_  & \new_Sorter100|13947_ ;
  assign \new_Sorter100|14047_  = \new_Sorter100|13946_  | \new_Sorter100|13947_ ;
  assign \new_Sorter100|14048_  = \new_Sorter100|13948_  & \new_Sorter100|13949_ ;
  assign \new_Sorter100|14049_  = \new_Sorter100|13948_  | \new_Sorter100|13949_ ;
  assign \new_Sorter100|14050_  = \new_Sorter100|13950_  & \new_Sorter100|13951_ ;
  assign \new_Sorter100|14051_  = \new_Sorter100|13950_  | \new_Sorter100|13951_ ;
  assign \new_Sorter100|14052_  = \new_Sorter100|13952_  & \new_Sorter100|13953_ ;
  assign \new_Sorter100|14053_  = \new_Sorter100|13952_  | \new_Sorter100|13953_ ;
  assign \new_Sorter100|14054_  = \new_Sorter100|13954_  & \new_Sorter100|13955_ ;
  assign \new_Sorter100|14055_  = \new_Sorter100|13954_  | \new_Sorter100|13955_ ;
  assign \new_Sorter100|14056_  = \new_Sorter100|13956_  & \new_Sorter100|13957_ ;
  assign \new_Sorter100|14057_  = \new_Sorter100|13956_  | \new_Sorter100|13957_ ;
  assign \new_Sorter100|14058_  = \new_Sorter100|13958_  & \new_Sorter100|13959_ ;
  assign \new_Sorter100|14059_  = \new_Sorter100|13958_  | \new_Sorter100|13959_ ;
  assign \new_Sorter100|14060_  = \new_Sorter100|13960_  & \new_Sorter100|13961_ ;
  assign \new_Sorter100|14061_  = \new_Sorter100|13960_  | \new_Sorter100|13961_ ;
  assign \new_Sorter100|14062_  = \new_Sorter100|13962_  & \new_Sorter100|13963_ ;
  assign \new_Sorter100|14063_  = \new_Sorter100|13962_  | \new_Sorter100|13963_ ;
  assign \new_Sorter100|14064_  = \new_Sorter100|13964_  & \new_Sorter100|13965_ ;
  assign \new_Sorter100|14065_  = \new_Sorter100|13964_  | \new_Sorter100|13965_ ;
  assign \new_Sorter100|14066_  = \new_Sorter100|13966_  & \new_Sorter100|13967_ ;
  assign \new_Sorter100|14067_  = \new_Sorter100|13966_  | \new_Sorter100|13967_ ;
  assign \new_Sorter100|14068_  = \new_Sorter100|13968_  & \new_Sorter100|13969_ ;
  assign \new_Sorter100|14069_  = \new_Sorter100|13968_  | \new_Sorter100|13969_ ;
  assign \new_Sorter100|14070_  = \new_Sorter100|13970_  & \new_Sorter100|13971_ ;
  assign \new_Sorter100|14071_  = \new_Sorter100|13970_  | \new_Sorter100|13971_ ;
  assign \new_Sorter100|14072_  = \new_Sorter100|13972_  & \new_Sorter100|13973_ ;
  assign \new_Sorter100|14073_  = \new_Sorter100|13972_  | \new_Sorter100|13973_ ;
  assign \new_Sorter100|14074_  = \new_Sorter100|13974_  & \new_Sorter100|13975_ ;
  assign \new_Sorter100|14075_  = \new_Sorter100|13974_  | \new_Sorter100|13975_ ;
  assign \new_Sorter100|14076_  = \new_Sorter100|13976_  & \new_Sorter100|13977_ ;
  assign \new_Sorter100|14077_  = \new_Sorter100|13976_  | \new_Sorter100|13977_ ;
  assign \new_Sorter100|14078_  = \new_Sorter100|13978_  & \new_Sorter100|13979_ ;
  assign \new_Sorter100|14079_  = \new_Sorter100|13978_  | \new_Sorter100|13979_ ;
  assign \new_Sorter100|14080_  = \new_Sorter100|13980_  & \new_Sorter100|13981_ ;
  assign \new_Sorter100|14081_  = \new_Sorter100|13980_  | \new_Sorter100|13981_ ;
  assign \new_Sorter100|14082_  = \new_Sorter100|13982_  & \new_Sorter100|13983_ ;
  assign \new_Sorter100|14083_  = \new_Sorter100|13982_  | \new_Sorter100|13983_ ;
  assign \new_Sorter100|14084_  = \new_Sorter100|13984_  & \new_Sorter100|13985_ ;
  assign \new_Sorter100|14085_  = \new_Sorter100|13984_  | \new_Sorter100|13985_ ;
  assign \new_Sorter100|14086_  = \new_Sorter100|13986_  & \new_Sorter100|13987_ ;
  assign \new_Sorter100|14087_  = \new_Sorter100|13986_  | \new_Sorter100|13987_ ;
  assign \new_Sorter100|14088_  = \new_Sorter100|13988_  & \new_Sorter100|13989_ ;
  assign \new_Sorter100|14089_  = \new_Sorter100|13988_  | \new_Sorter100|13989_ ;
  assign \new_Sorter100|14090_  = \new_Sorter100|13990_  & \new_Sorter100|13991_ ;
  assign \new_Sorter100|14091_  = \new_Sorter100|13990_  | \new_Sorter100|13991_ ;
  assign \new_Sorter100|14092_  = \new_Sorter100|13992_  & \new_Sorter100|13993_ ;
  assign \new_Sorter100|14093_  = \new_Sorter100|13992_  | \new_Sorter100|13993_ ;
  assign \new_Sorter100|14094_  = \new_Sorter100|13994_  & \new_Sorter100|13995_ ;
  assign \new_Sorter100|14095_  = \new_Sorter100|13994_  | \new_Sorter100|13995_ ;
  assign \new_Sorter100|14096_  = \new_Sorter100|13996_  & \new_Sorter100|13997_ ;
  assign \new_Sorter100|14097_  = \new_Sorter100|13996_  | \new_Sorter100|13997_ ;
  assign \new_Sorter100|14098_  = \new_Sorter100|13998_  & \new_Sorter100|13999_ ;
  assign \new_Sorter100|14099_  = \new_Sorter100|13998_  | \new_Sorter100|13999_ ;
  assign \new_Sorter100|14100_  = \new_Sorter100|14000_ ;
  assign \new_Sorter100|14199_  = \new_Sorter100|14099_ ;
  assign \new_Sorter100|14101_  = \new_Sorter100|14001_  & \new_Sorter100|14002_ ;
  assign \new_Sorter100|14102_  = \new_Sorter100|14001_  | \new_Sorter100|14002_ ;
  assign \new_Sorter100|14103_  = \new_Sorter100|14003_  & \new_Sorter100|14004_ ;
  assign \new_Sorter100|14104_  = \new_Sorter100|14003_  | \new_Sorter100|14004_ ;
  assign \new_Sorter100|14105_  = \new_Sorter100|14005_  & \new_Sorter100|14006_ ;
  assign \new_Sorter100|14106_  = \new_Sorter100|14005_  | \new_Sorter100|14006_ ;
  assign \new_Sorter100|14107_  = \new_Sorter100|14007_  & \new_Sorter100|14008_ ;
  assign \new_Sorter100|14108_  = \new_Sorter100|14007_  | \new_Sorter100|14008_ ;
  assign \new_Sorter100|14109_  = \new_Sorter100|14009_  & \new_Sorter100|14010_ ;
  assign \new_Sorter100|14110_  = \new_Sorter100|14009_  | \new_Sorter100|14010_ ;
  assign \new_Sorter100|14111_  = \new_Sorter100|14011_  & \new_Sorter100|14012_ ;
  assign \new_Sorter100|14112_  = \new_Sorter100|14011_  | \new_Sorter100|14012_ ;
  assign \new_Sorter100|14113_  = \new_Sorter100|14013_  & \new_Sorter100|14014_ ;
  assign \new_Sorter100|14114_  = \new_Sorter100|14013_  | \new_Sorter100|14014_ ;
  assign \new_Sorter100|14115_  = \new_Sorter100|14015_  & \new_Sorter100|14016_ ;
  assign \new_Sorter100|14116_  = \new_Sorter100|14015_  | \new_Sorter100|14016_ ;
  assign \new_Sorter100|14117_  = \new_Sorter100|14017_  & \new_Sorter100|14018_ ;
  assign \new_Sorter100|14118_  = \new_Sorter100|14017_  | \new_Sorter100|14018_ ;
  assign \new_Sorter100|14119_  = \new_Sorter100|14019_  & \new_Sorter100|14020_ ;
  assign \new_Sorter100|14120_  = \new_Sorter100|14019_  | \new_Sorter100|14020_ ;
  assign \new_Sorter100|14121_  = \new_Sorter100|14021_  & \new_Sorter100|14022_ ;
  assign \new_Sorter100|14122_  = \new_Sorter100|14021_  | \new_Sorter100|14022_ ;
  assign \new_Sorter100|14123_  = \new_Sorter100|14023_  & \new_Sorter100|14024_ ;
  assign \new_Sorter100|14124_  = \new_Sorter100|14023_  | \new_Sorter100|14024_ ;
  assign \new_Sorter100|14125_  = \new_Sorter100|14025_  & \new_Sorter100|14026_ ;
  assign \new_Sorter100|14126_  = \new_Sorter100|14025_  | \new_Sorter100|14026_ ;
  assign \new_Sorter100|14127_  = \new_Sorter100|14027_  & \new_Sorter100|14028_ ;
  assign \new_Sorter100|14128_  = \new_Sorter100|14027_  | \new_Sorter100|14028_ ;
  assign \new_Sorter100|14129_  = \new_Sorter100|14029_  & \new_Sorter100|14030_ ;
  assign \new_Sorter100|14130_  = \new_Sorter100|14029_  | \new_Sorter100|14030_ ;
  assign \new_Sorter100|14131_  = \new_Sorter100|14031_  & \new_Sorter100|14032_ ;
  assign \new_Sorter100|14132_  = \new_Sorter100|14031_  | \new_Sorter100|14032_ ;
  assign \new_Sorter100|14133_  = \new_Sorter100|14033_  & \new_Sorter100|14034_ ;
  assign \new_Sorter100|14134_  = \new_Sorter100|14033_  | \new_Sorter100|14034_ ;
  assign \new_Sorter100|14135_  = \new_Sorter100|14035_  & \new_Sorter100|14036_ ;
  assign \new_Sorter100|14136_  = \new_Sorter100|14035_  | \new_Sorter100|14036_ ;
  assign \new_Sorter100|14137_  = \new_Sorter100|14037_  & \new_Sorter100|14038_ ;
  assign \new_Sorter100|14138_  = \new_Sorter100|14037_  | \new_Sorter100|14038_ ;
  assign \new_Sorter100|14139_  = \new_Sorter100|14039_  & \new_Sorter100|14040_ ;
  assign \new_Sorter100|14140_  = \new_Sorter100|14039_  | \new_Sorter100|14040_ ;
  assign \new_Sorter100|14141_  = \new_Sorter100|14041_  & \new_Sorter100|14042_ ;
  assign \new_Sorter100|14142_  = \new_Sorter100|14041_  | \new_Sorter100|14042_ ;
  assign \new_Sorter100|14143_  = \new_Sorter100|14043_  & \new_Sorter100|14044_ ;
  assign \new_Sorter100|14144_  = \new_Sorter100|14043_  | \new_Sorter100|14044_ ;
  assign \new_Sorter100|14145_  = \new_Sorter100|14045_  & \new_Sorter100|14046_ ;
  assign \new_Sorter100|14146_  = \new_Sorter100|14045_  | \new_Sorter100|14046_ ;
  assign \new_Sorter100|14147_  = \new_Sorter100|14047_  & \new_Sorter100|14048_ ;
  assign \new_Sorter100|14148_  = \new_Sorter100|14047_  | \new_Sorter100|14048_ ;
  assign \new_Sorter100|14149_  = \new_Sorter100|14049_  & \new_Sorter100|14050_ ;
  assign \new_Sorter100|14150_  = \new_Sorter100|14049_  | \new_Sorter100|14050_ ;
  assign \new_Sorter100|14151_  = \new_Sorter100|14051_  & \new_Sorter100|14052_ ;
  assign \new_Sorter100|14152_  = \new_Sorter100|14051_  | \new_Sorter100|14052_ ;
  assign \new_Sorter100|14153_  = \new_Sorter100|14053_  & \new_Sorter100|14054_ ;
  assign \new_Sorter100|14154_  = \new_Sorter100|14053_  | \new_Sorter100|14054_ ;
  assign \new_Sorter100|14155_  = \new_Sorter100|14055_  & \new_Sorter100|14056_ ;
  assign \new_Sorter100|14156_  = \new_Sorter100|14055_  | \new_Sorter100|14056_ ;
  assign \new_Sorter100|14157_  = \new_Sorter100|14057_  & \new_Sorter100|14058_ ;
  assign \new_Sorter100|14158_  = \new_Sorter100|14057_  | \new_Sorter100|14058_ ;
  assign \new_Sorter100|14159_  = \new_Sorter100|14059_  & \new_Sorter100|14060_ ;
  assign \new_Sorter100|14160_  = \new_Sorter100|14059_  | \new_Sorter100|14060_ ;
  assign \new_Sorter100|14161_  = \new_Sorter100|14061_  & \new_Sorter100|14062_ ;
  assign \new_Sorter100|14162_  = \new_Sorter100|14061_  | \new_Sorter100|14062_ ;
  assign \new_Sorter100|14163_  = \new_Sorter100|14063_  & \new_Sorter100|14064_ ;
  assign \new_Sorter100|14164_  = \new_Sorter100|14063_  | \new_Sorter100|14064_ ;
  assign \new_Sorter100|14165_  = \new_Sorter100|14065_  & \new_Sorter100|14066_ ;
  assign \new_Sorter100|14166_  = \new_Sorter100|14065_  | \new_Sorter100|14066_ ;
  assign \new_Sorter100|14167_  = \new_Sorter100|14067_  & \new_Sorter100|14068_ ;
  assign \new_Sorter100|14168_  = \new_Sorter100|14067_  | \new_Sorter100|14068_ ;
  assign \new_Sorter100|14169_  = \new_Sorter100|14069_  & \new_Sorter100|14070_ ;
  assign \new_Sorter100|14170_  = \new_Sorter100|14069_  | \new_Sorter100|14070_ ;
  assign \new_Sorter100|14171_  = \new_Sorter100|14071_  & \new_Sorter100|14072_ ;
  assign \new_Sorter100|14172_  = \new_Sorter100|14071_  | \new_Sorter100|14072_ ;
  assign \new_Sorter100|14173_  = \new_Sorter100|14073_  & \new_Sorter100|14074_ ;
  assign \new_Sorter100|14174_  = \new_Sorter100|14073_  | \new_Sorter100|14074_ ;
  assign \new_Sorter100|14175_  = \new_Sorter100|14075_  & \new_Sorter100|14076_ ;
  assign \new_Sorter100|14176_  = \new_Sorter100|14075_  | \new_Sorter100|14076_ ;
  assign \new_Sorter100|14177_  = \new_Sorter100|14077_  & \new_Sorter100|14078_ ;
  assign \new_Sorter100|14178_  = \new_Sorter100|14077_  | \new_Sorter100|14078_ ;
  assign \new_Sorter100|14179_  = \new_Sorter100|14079_  & \new_Sorter100|14080_ ;
  assign \new_Sorter100|14180_  = \new_Sorter100|14079_  | \new_Sorter100|14080_ ;
  assign \new_Sorter100|14181_  = \new_Sorter100|14081_  & \new_Sorter100|14082_ ;
  assign \new_Sorter100|14182_  = \new_Sorter100|14081_  | \new_Sorter100|14082_ ;
  assign \new_Sorter100|14183_  = \new_Sorter100|14083_  & \new_Sorter100|14084_ ;
  assign \new_Sorter100|14184_  = \new_Sorter100|14083_  | \new_Sorter100|14084_ ;
  assign \new_Sorter100|14185_  = \new_Sorter100|14085_  & \new_Sorter100|14086_ ;
  assign \new_Sorter100|14186_  = \new_Sorter100|14085_  | \new_Sorter100|14086_ ;
  assign \new_Sorter100|14187_  = \new_Sorter100|14087_  & \new_Sorter100|14088_ ;
  assign \new_Sorter100|14188_  = \new_Sorter100|14087_  | \new_Sorter100|14088_ ;
  assign \new_Sorter100|14189_  = \new_Sorter100|14089_  & \new_Sorter100|14090_ ;
  assign \new_Sorter100|14190_  = \new_Sorter100|14089_  | \new_Sorter100|14090_ ;
  assign \new_Sorter100|14191_  = \new_Sorter100|14091_  & \new_Sorter100|14092_ ;
  assign \new_Sorter100|14192_  = \new_Sorter100|14091_  | \new_Sorter100|14092_ ;
  assign \new_Sorter100|14193_  = \new_Sorter100|14093_  & \new_Sorter100|14094_ ;
  assign \new_Sorter100|14194_  = \new_Sorter100|14093_  | \new_Sorter100|14094_ ;
  assign \new_Sorter100|14195_  = \new_Sorter100|14095_  & \new_Sorter100|14096_ ;
  assign \new_Sorter100|14196_  = \new_Sorter100|14095_  | \new_Sorter100|14096_ ;
  assign \new_Sorter100|14197_  = \new_Sorter100|14097_  & \new_Sorter100|14098_ ;
  assign \new_Sorter100|14198_  = \new_Sorter100|14097_  | \new_Sorter100|14098_ ;
  assign \new_Sorter100|14200_  = \new_Sorter100|14100_  & \new_Sorter100|14101_ ;
  assign \new_Sorter100|14201_  = \new_Sorter100|14100_  | \new_Sorter100|14101_ ;
  assign \new_Sorter100|14202_  = \new_Sorter100|14102_  & \new_Sorter100|14103_ ;
  assign \new_Sorter100|14203_  = \new_Sorter100|14102_  | \new_Sorter100|14103_ ;
  assign \new_Sorter100|14204_  = \new_Sorter100|14104_  & \new_Sorter100|14105_ ;
  assign \new_Sorter100|14205_  = \new_Sorter100|14104_  | \new_Sorter100|14105_ ;
  assign \new_Sorter100|14206_  = \new_Sorter100|14106_  & \new_Sorter100|14107_ ;
  assign \new_Sorter100|14207_  = \new_Sorter100|14106_  | \new_Sorter100|14107_ ;
  assign \new_Sorter100|14208_  = \new_Sorter100|14108_  & \new_Sorter100|14109_ ;
  assign \new_Sorter100|14209_  = \new_Sorter100|14108_  | \new_Sorter100|14109_ ;
  assign \new_Sorter100|14210_  = \new_Sorter100|14110_  & \new_Sorter100|14111_ ;
  assign \new_Sorter100|14211_  = \new_Sorter100|14110_  | \new_Sorter100|14111_ ;
  assign \new_Sorter100|14212_  = \new_Sorter100|14112_  & \new_Sorter100|14113_ ;
  assign \new_Sorter100|14213_  = \new_Sorter100|14112_  | \new_Sorter100|14113_ ;
  assign \new_Sorter100|14214_  = \new_Sorter100|14114_  & \new_Sorter100|14115_ ;
  assign \new_Sorter100|14215_  = \new_Sorter100|14114_  | \new_Sorter100|14115_ ;
  assign \new_Sorter100|14216_  = \new_Sorter100|14116_  & \new_Sorter100|14117_ ;
  assign \new_Sorter100|14217_  = \new_Sorter100|14116_  | \new_Sorter100|14117_ ;
  assign \new_Sorter100|14218_  = \new_Sorter100|14118_  & \new_Sorter100|14119_ ;
  assign \new_Sorter100|14219_  = \new_Sorter100|14118_  | \new_Sorter100|14119_ ;
  assign \new_Sorter100|14220_  = \new_Sorter100|14120_  & \new_Sorter100|14121_ ;
  assign \new_Sorter100|14221_  = \new_Sorter100|14120_  | \new_Sorter100|14121_ ;
  assign \new_Sorter100|14222_  = \new_Sorter100|14122_  & \new_Sorter100|14123_ ;
  assign \new_Sorter100|14223_  = \new_Sorter100|14122_  | \new_Sorter100|14123_ ;
  assign \new_Sorter100|14224_  = \new_Sorter100|14124_  & \new_Sorter100|14125_ ;
  assign \new_Sorter100|14225_  = \new_Sorter100|14124_  | \new_Sorter100|14125_ ;
  assign \new_Sorter100|14226_  = \new_Sorter100|14126_  & \new_Sorter100|14127_ ;
  assign \new_Sorter100|14227_  = \new_Sorter100|14126_  | \new_Sorter100|14127_ ;
  assign \new_Sorter100|14228_  = \new_Sorter100|14128_  & \new_Sorter100|14129_ ;
  assign \new_Sorter100|14229_  = \new_Sorter100|14128_  | \new_Sorter100|14129_ ;
  assign \new_Sorter100|14230_  = \new_Sorter100|14130_  & \new_Sorter100|14131_ ;
  assign \new_Sorter100|14231_  = \new_Sorter100|14130_  | \new_Sorter100|14131_ ;
  assign \new_Sorter100|14232_  = \new_Sorter100|14132_  & \new_Sorter100|14133_ ;
  assign \new_Sorter100|14233_  = \new_Sorter100|14132_  | \new_Sorter100|14133_ ;
  assign \new_Sorter100|14234_  = \new_Sorter100|14134_  & \new_Sorter100|14135_ ;
  assign \new_Sorter100|14235_  = \new_Sorter100|14134_  | \new_Sorter100|14135_ ;
  assign \new_Sorter100|14236_  = \new_Sorter100|14136_  & \new_Sorter100|14137_ ;
  assign \new_Sorter100|14237_  = \new_Sorter100|14136_  | \new_Sorter100|14137_ ;
  assign \new_Sorter100|14238_  = \new_Sorter100|14138_  & \new_Sorter100|14139_ ;
  assign \new_Sorter100|14239_  = \new_Sorter100|14138_  | \new_Sorter100|14139_ ;
  assign \new_Sorter100|14240_  = \new_Sorter100|14140_  & \new_Sorter100|14141_ ;
  assign \new_Sorter100|14241_  = \new_Sorter100|14140_  | \new_Sorter100|14141_ ;
  assign \new_Sorter100|14242_  = \new_Sorter100|14142_  & \new_Sorter100|14143_ ;
  assign \new_Sorter100|14243_  = \new_Sorter100|14142_  | \new_Sorter100|14143_ ;
  assign \new_Sorter100|14244_  = \new_Sorter100|14144_  & \new_Sorter100|14145_ ;
  assign \new_Sorter100|14245_  = \new_Sorter100|14144_  | \new_Sorter100|14145_ ;
  assign \new_Sorter100|14246_  = \new_Sorter100|14146_  & \new_Sorter100|14147_ ;
  assign \new_Sorter100|14247_  = \new_Sorter100|14146_  | \new_Sorter100|14147_ ;
  assign \new_Sorter100|14248_  = \new_Sorter100|14148_  & \new_Sorter100|14149_ ;
  assign \new_Sorter100|14249_  = \new_Sorter100|14148_  | \new_Sorter100|14149_ ;
  assign \new_Sorter100|14250_  = \new_Sorter100|14150_  & \new_Sorter100|14151_ ;
  assign \new_Sorter100|14251_  = \new_Sorter100|14150_  | \new_Sorter100|14151_ ;
  assign \new_Sorter100|14252_  = \new_Sorter100|14152_  & \new_Sorter100|14153_ ;
  assign \new_Sorter100|14253_  = \new_Sorter100|14152_  | \new_Sorter100|14153_ ;
  assign \new_Sorter100|14254_  = \new_Sorter100|14154_  & \new_Sorter100|14155_ ;
  assign \new_Sorter100|14255_  = \new_Sorter100|14154_  | \new_Sorter100|14155_ ;
  assign \new_Sorter100|14256_  = \new_Sorter100|14156_  & \new_Sorter100|14157_ ;
  assign \new_Sorter100|14257_  = \new_Sorter100|14156_  | \new_Sorter100|14157_ ;
  assign \new_Sorter100|14258_  = \new_Sorter100|14158_  & \new_Sorter100|14159_ ;
  assign \new_Sorter100|14259_  = \new_Sorter100|14158_  | \new_Sorter100|14159_ ;
  assign \new_Sorter100|14260_  = \new_Sorter100|14160_  & \new_Sorter100|14161_ ;
  assign \new_Sorter100|14261_  = \new_Sorter100|14160_  | \new_Sorter100|14161_ ;
  assign \new_Sorter100|14262_  = \new_Sorter100|14162_  & \new_Sorter100|14163_ ;
  assign \new_Sorter100|14263_  = \new_Sorter100|14162_  | \new_Sorter100|14163_ ;
  assign \new_Sorter100|14264_  = \new_Sorter100|14164_  & \new_Sorter100|14165_ ;
  assign \new_Sorter100|14265_  = \new_Sorter100|14164_  | \new_Sorter100|14165_ ;
  assign \new_Sorter100|14266_  = \new_Sorter100|14166_  & \new_Sorter100|14167_ ;
  assign \new_Sorter100|14267_  = \new_Sorter100|14166_  | \new_Sorter100|14167_ ;
  assign \new_Sorter100|14268_  = \new_Sorter100|14168_  & \new_Sorter100|14169_ ;
  assign \new_Sorter100|14269_  = \new_Sorter100|14168_  | \new_Sorter100|14169_ ;
  assign \new_Sorter100|14270_  = \new_Sorter100|14170_  & \new_Sorter100|14171_ ;
  assign \new_Sorter100|14271_  = \new_Sorter100|14170_  | \new_Sorter100|14171_ ;
  assign \new_Sorter100|14272_  = \new_Sorter100|14172_  & \new_Sorter100|14173_ ;
  assign \new_Sorter100|14273_  = \new_Sorter100|14172_  | \new_Sorter100|14173_ ;
  assign \new_Sorter100|14274_  = \new_Sorter100|14174_  & \new_Sorter100|14175_ ;
  assign \new_Sorter100|14275_  = \new_Sorter100|14174_  | \new_Sorter100|14175_ ;
  assign \new_Sorter100|14276_  = \new_Sorter100|14176_  & \new_Sorter100|14177_ ;
  assign \new_Sorter100|14277_  = \new_Sorter100|14176_  | \new_Sorter100|14177_ ;
  assign \new_Sorter100|14278_  = \new_Sorter100|14178_  & \new_Sorter100|14179_ ;
  assign \new_Sorter100|14279_  = \new_Sorter100|14178_  | \new_Sorter100|14179_ ;
  assign \new_Sorter100|14280_  = \new_Sorter100|14180_  & \new_Sorter100|14181_ ;
  assign \new_Sorter100|14281_  = \new_Sorter100|14180_  | \new_Sorter100|14181_ ;
  assign \new_Sorter100|14282_  = \new_Sorter100|14182_  & \new_Sorter100|14183_ ;
  assign \new_Sorter100|14283_  = \new_Sorter100|14182_  | \new_Sorter100|14183_ ;
  assign \new_Sorter100|14284_  = \new_Sorter100|14184_  & \new_Sorter100|14185_ ;
  assign \new_Sorter100|14285_  = \new_Sorter100|14184_  | \new_Sorter100|14185_ ;
  assign \new_Sorter100|14286_  = \new_Sorter100|14186_  & \new_Sorter100|14187_ ;
  assign \new_Sorter100|14287_  = \new_Sorter100|14186_  | \new_Sorter100|14187_ ;
  assign \new_Sorter100|14288_  = \new_Sorter100|14188_  & \new_Sorter100|14189_ ;
  assign \new_Sorter100|14289_  = \new_Sorter100|14188_  | \new_Sorter100|14189_ ;
  assign \new_Sorter100|14290_  = \new_Sorter100|14190_  & \new_Sorter100|14191_ ;
  assign \new_Sorter100|14291_  = \new_Sorter100|14190_  | \new_Sorter100|14191_ ;
  assign \new_Sorter100|14292_  = \new_Sorter100|14192_  & \new_Sorter100|14193_ ;
  assign \new_Sorter100|14293_  = \new_Sorter100|14192_  | \new_Sorter100|14193_ ;
  assign \new_Sorter100|14294_  = \new_Sorter100|14194_  & \new_Sorter100|14195_ ;
  assign \new_Sorter100|14295_  = \new_Sorter100|14194_  | \new_Sorter100|14195_ ;
  assign \new_Sorter100|14296_  = \new_Sorter100|14196_  & \new_Sorter100|14197_ ;
  assign \new_Sorter100|14297_  = \new_Sorter100|14196_  | \new_Sorter100|14197_ ;
  assign \new_Sorter100|14298_  = \new_Sorter100|14198_  & \new_Sorter100|14199_ ;
  assign \new_Sorter100|14299_  = \new_Sorter100|14198_  | \new_Sorter100|14199_ ;
  assign \new_Sorter100|14300_  = \new_Sorter100|14200_ ;
  assign \new_Sorter100|14399_  = \new_Sorter100|14299_ ;
  assign \new_Sorter100|14301_  = \new_Sorter100|14201_  & \new_Sorter100|14202_ ;
  assign \new_Sorter100|14302_  = \new_Sorter100|14201_  | \new_Sorter100|14202_ ;
  assign \new_Sorter100|14303_  = \new_Sorter100|14203_  & \new_Sorter100|14204_ ;
  assign \new_Sorter100|14304_  = \new_Sorter100|14203_  | \new_Sorter100|14204_ ;
  assign \new_Sorter100|14305_  = \new_Sorter100|14205_  & \new_Sorter100|14206_ ;
  assign \new_Sorter100|14306_  = \new_Sorter100|14205_  | \new_Sorter100|14206_ ;
  assign \new_Sorter100|14307_  = \new_Sorter100|14207_  & \new_Sorter100|14208_ ;
  assign \new_Sorter100|14308_  = \new_Sorter100|14207_  | \new_Sorter100|14208_ ;
  assign \new_Sorter100|14309_  = \new_Sorter100|14209_  & \new_Sorter100|14210_ ;
  assign \new_Sorter100|14310_  = \new_Sorter100|14209_  | \new_Sorter100|14210_ ;
  assign \new_Sorter100|14311_  = \new_Sorter100|14211_  & \new_Sorter100|14212_ ;
  assign \new_Sorter100|14312_  = \new_Sorter100|14211_  | \new_Sorter100|14212_ ;
  assign \new_Sorter100|14313_  = \new_Sorter100|14213_  & \new_Sorter100|14214_ ;
  assign \new_Sorter100|14314_  = \new_Sorter100|14213_  | \new_Sorter100|14214_ ;
  assign \new_Sorter100|14315_  = \new_Sorter100|14215_  & \new_Sorter100|14216_ ;
  assign \new_Sorter100|14316_  = \new_Sorter100|14215_  | \new_Sorter100|14216_ ;
  assign \new_Sorter100|14317_  = \new_Sorter100|14217_  & \new_Sorter100|14218_ ;
  assign \new_Sorter100|14318_  = \new_Sorter100|14217_  | \new_Sorter100|14218_ ;
  assign \new_Sorter100|14319_  = \new_Sorter100|14219_  & \new_Sorter100|14220_ ;
  assign \new_Sorter100|14320_  = \new_Sorter100|14219_  | \new_Sorter100|14220_ ;
  assign \new_Sorter100|14321_  = \new_Sorter100|14221_  & \new_Sorter100|14222_ ;
  assign \new_Sorter100|14322_  = \new_Sorter100|14221_  | \new_Sorter100|14222_ ;
  assign \new_Sorter100|14323_  = \new_Sorter100|14223_  & \new_Sorter100|14224_ ;
  assign \new_Sorter100|14324_  = \new_Sorter100|14223_  | \new_Sorter100|14224_ ;
  assign \new_Sorter100|14325_  = \new_Sorter100|14225_  & \new_Sorter100|14226_ ;
  assign \new_Sorter100|14326_  = \new_Sorter100|14225_  | \new_Sorter100|14226_ ;
  assign \new_Sorter100|14327_  = \new_Sorter100|14227_  & \new_Sorter100|14228_ ;
  assign \new_Sorter100|14328_  = \new_Sorter100|14227_  | \new_Sorter100|14228_ ;
  assign \new_Sorter100|14329_  = \new_Sorter100|14229_  & \new_Sorter100|14230_ ;
  assign \new_Sorter100|14330_  = \new_Sorter100|14229_  | \new_Sorter100|14230_ ;
  assign \new_Sorter100|14331_  = \new_Sorter100|14231_  & \new_Sorter100|14232_ ;
  assign \new_Sorter100|14332_  = \new_Sorter100|14231_  | \new_Sorter100|14232_ ;
  assign \new_Sorter100|14333_  = \new_Sorter100|14233_  & \new_Sorter100|14234_ ;
  assign \new_Sorter100|14334_  = \new_Sorter100|14233_  | \new_Sorter100|14234_ ;
  assign \new_Sorter100|14335_  = \new_Sorter100|14235_  & \new_Sorter100|14236_ ;
  assign \new_Sorter100|14336_  = \new_Sorter100|14235_  | \new_Sorter100|14236_ ;
  assign \new_Sorter100|14337_  = \new_Sorter100|14237_  & \new_Sorter100|14238_ ;
  assign \new_Sorter100|14338_  = \new_Sorter100|14237_  | \new_Sorter100|14238_ ;
  assign \new_Sorter100|14339_  = \new_Sorter100|14239_  & \new_Sorter100|14240_ ;
  assign \new_Sorter100|14340_  = \new_Sorter100|14239_  | \new_Sorter100|14240_ ;
  assign \new_Sorter100|14341_  = \new_Sorter100|14241_  & \new_Sorter100|14242_ ;
  assign \new_Sorter100|14342_  = \new_Sorter100|14241_  | \new_Sorter100|14242_ ;
  assign \new_Sorter100|14343_  = \new_Sorter100|14243_  & \new_Sorter100|14244_ ;
  assign \new_Sorter100|14344_  = \new_Sorter100|14243_  | \new_Sorter100|14244_ ;
  assign \new_Sorter100|14345_  = \new_Sorter100|14245_  & \new_Sorter100|14246_ ;
  assign \new_Sorter100|14346_  = \new_Sorter100|14245_  | \new_Sorter100|14246_ ;
  assign \new_Sorter100|14347_  = \new_Sorter100|14247_  & \new_Sorter100|14248_ ;
  assign \new_Sorter100|14348_  = \new_Sorter100|14247_  | \new_Sorter100|14248_ ;
  assign \new_Sorter100|14349_  = \new_Sorter100|14249_  & \new_Sorter100|14250_ ;
  assign \new_Sorter100|14350_  = \new_Sorter100|14249_  | \new_Sorter100|14250_ ;
  assign \new_Sorter100|14351_  = \new_Sorter100|14251_  & \new_Sorter100|14252_ ;
  assign \new_Sorter100|14352_  = \new_Sorter100|14251_  | \new_Sorter100|14252_ ;
  assign \new_Sorter100|14353_  = \new_Sorter100|14253_  & \new_Sorter100|14254_ ;
  assign \new_Sorter100|14354_  = \new_Sorter100|14253_  | \new_Sorter100|14254_ ;
  assign \new_Sorter100|14355_  = \new_Sorter100|14255_  & \new_Sorter100|14256_ ;
  assign \new_Sorter100|14356_  = \new_Sorter100|14255_  | \new_Sorter100|14256_ ;
  assign \new_Sorter100|14357_  = \new_Sorter100|14257_  & \new_Sorter100|14258_ ;
  assign \new_Sorter100|14358_  = \new_Sorter100|14257_  | \new_Sorter100|14258_ ;
  assign \new_Sorter100|14359_  = \new_Sorter100|14259_  & \new_Sorter100|14260_ ;
  assign \new_Sorter100|14360_  = \new_Sorter100|14259_  | \new_Sorter100|14260_ ;
  assign \new_Sorter100|14361_  = \new_Sorter100|14261_  & \new_Sorter100|14262_ ;
  assign \new_Sorter100|14362_  = \new_Sorter100|14261_  | \new_Sorter100|14262_ ;
  assign \new_Sorter100|14363_  = \new_Sorter100|14263_  & \new_Sorter100|14264_ ;
  assign \new_Sorter100|14364_  = \new_Sorter100|14263_  | \new_Sorter100|14264_ ;
  assign \new_Sorter100|14365_  = \new_Sorter100|14265_  & \new_Sorter100|14266_ ;
  assign \new_Sorter100|14366_  = \new_Sorter100|14265_  | \new_Sorter100|14266_ ;
  assign \new_Sorter100|14367_  = \new_Sorter100|14267_  & \new_Sorter100|14268_ ;
  assign \new_Sorter100|14368_  = \new_Sorter100|14267_  | \new_Sorter100|14268_ ;
  assign \new_Sorter100|14369_  = \new_Sorter100|14269_  & \new_Sorter100|14270_ ;
  assign \new_Sorter100|14370_  = \new_Sorter100|14269_  | \new_Sorter100|14270_ ;
  assign \new_Sorter100|14371_  = \new_Sorter100|14271_  & \new_Sorter100|14272_ ;
  assign \new_Sorter100|14372_  = \new_Sorter100|14271_  | \new_Sorter100|14272_ ;
  assign \new_Sorter100|14373_  = \new_Sorter100|14273_  & \new_Sorter100|14274_ ;
  assign \new_Sorter100|14374_  = \new_Sorter100|14273_  | \new_Sorter100|14274_ ;
  assign \new_Sorter100|14375_  = \new_Sorter100|14275_  & \new_Sorter100|14276_ ;
  assign \new_Sorter100|14376_  = \new_Sorter100|14275_  | \new_Sorter100|14276_ ;
  assign \new_Sorter100|14377_  = \new_Sorter100|14277_  & \new_Sorter100|14278_ ;
  assign \new_Sorter100|14378_  = \new_Sorter100|14277_  | \new_Sorter100|14278_ ;
  assign \new_Sorter100|14379_  = \new_Sorter100|14279_  & \new_Sorter100|14280_ ;
  assign \new_Sorter100|14380_  = \new_Sorter100|14279_  | \new_Sorter100|14280_ ;
  assign \new_Sorter100|14381_  = \new_Sorter100|14281_  & \new_Sorter100|14282_ ;
  assign \new_Sorter100|14382_  = \new_Sorter100|14281_  | \new_Sorter100|14282_ ;
  assign \new_Sorter100|14383_  = \new_Sorter100|14283_  & \new_Sorter100|14284_ ;
  assign \new_Sorter100|14384_  = \new_Sorter100|14283_  | \new_Sorter100|14284_ ;
  assign \new_Sorter100|14385_  = \new_Sorter100|14285_  & \new_Sorter100|14286_ ;
  assign \new_Sorter100|14386_  = \new_Sorter100|14285_  | \new_Sorter100|14286_ ;
  assign \new_Sorter100|14387_  = \new_Sorter100|14287_  & \new_Sorter100|14288_ ;
  assign \new_Sorter100|14388_  = \new_Sorter100|14287_  | \new_Sorter100|14288_ ;
  assign \new_Sorter100|14389_  = \new_Sorter100|14289_  & \new_Sorter100|14290_ ;
  assign \new_Sorter100|14390_  = \new_Sorter100|14289_  | \new_Sorter100|14290_ ;
  assign \new_Sorter100|14391_  = \new_Sorter100|14291_  & \new_Sorter100|14292_ ;
  assign \new_Sorter100|14392_  = \new_Sorter100|14291_  | \new_Sorter100|14292_ ;
  assign \new_Sorter100|14393_  = \new_Sorter100|14293_  & \new_Sorter100|14294_ ;
  assign \new_Sorter100|14394_  = \new_Sorter100|14293_  | \new_Sorter100|14294_ ;
  assign \new_Sorter100|14395_  = \new_Sorter100|14295_  & \new_Sorter100|14296_ ;
  assign \new_Sorter100|14396_  = \new_Sorter100|14295_  | \new_Sorter100|14296_ ;
  assign \new_Sorter100|14397_  = \new_Sorter100|14297_  & \new_Sorter100|14298_ ;
  assign \new_Sorter100|14398_  = \new_Sorter100|14297_  | \new_Sorter100|14298_ ;
  assign \new_Sorter100|14400_  = \new_Sorter100|14300_  & \new_Sorter100|14301_ ;
  assign \new_Sorter100|14401_  = \new_Sorter100|14300_  | \new_Sorter100|14301_ ;
  assign \new_Sorter100|14402_  = \new_Sorter100|14302_  & \new_Sorter100|14303_ ;
  assign \new_Sorter100|14403_  = \new_Sorter100|14302_  | \new_Sorter100|14303_ ;
  assign \new_Sorter100|14404_  = \new_Sorter100|14304_  & \new_Sorter100|14305_ ;
  assign \new_Sorter100|14405_  = \new_Sorter100|14304_  | \new_Sorter100|14305_ ;
  assign \new_Sorter100|14406_  = \new_Sorter100|14306_  & \new_Sorter100|14307_ ;
  assign \new_Sorter100|14407_  = \new_Sorter100|14306_  | \new_Sorter100|14307_ ;
  assign \new_Sorter100|14408_  = \new_Sorter100|14308_  & \new_Sorter100|14309_ ;
  assign \new_Sorter100|14409_  = \new_Sorter100|14308_  | \new_Sorter100|14309_ ;
  assign \new_Sorter100|14410_  = \new_Sorter100|14310_  & \new_Sorter100|14311_ ;
  assign \new_Sorter100|14411_  = \new_Sorter100|14310_  | \new_Sorter100|14311_ ;
  assign \new_Sorter100|14412_  = \new_Sorter100|14312_  & \new_Sorter100|14313_ ;
  assign \new_Sorter100|14413_  = \new_Sorter100|14312_  | \new_Sorter100|14313_ ;
  assign \new_Sorter100|14414_  = \new_Sorter100|14314_  & \new_Sorter100|14315_ ;
  assign \new_Sorter100|14415_  = \new_Sorter100|14314_  | \new_Sorter100|14315_ ;
  assign \new_Sorter100|14416_  = \new_Sorter100|14316_  & \new_Sorter100|14317_ ;
  assign \new_Sorter100|14417_  = \new_Sorter100|14316_  | \new_Sorter100|14317_ ;
  assign \new_Sorter100|14418_  = \new_Sorter100|14318_  & \new_Sorter100|14319_ ;
  assign \new_Sorter100|14419_  = \new_Sorter100|14318_  | \new_Sorter100|14319_ ;
  assign \new_Sorter100|14420_  = \new_Sorter100|14320_  & \new_Sorter100|14321_ ;
  assign \new_Sorter100|14421_  = \new_Sorter100|14320_  | \new_Sorter100|14321_ ;
  assign \new_Sorter100|14422_  = \new_Sorter100|14322_  & \new_Sorter100|14323_ ;
  assign \new_Sorter100|14423_  = \new_Sorter100|14322_  | \new_Sorter100|14323_ ;
  assign \new_Sorter100|14424_  = \new_Sorter100|14324_  & \new_Sorter100|14325_ ;
  assign \new_Sorter100|14425_  = \new_Sorter100|14324_  | \new_Sorter100|14325_ ;
  assign \new_Sorter100|14426_  = \new_Sorter100|14326_  & \new_Sorter100|14327_ ;
  assign \new_Sorter100|14427_  = \new_Sorter100|14326_  | \new_Sorter100|14327_ ;
  assign \new_Sorter100|14428_  = \new_Sorter100|14328_  & \new_Sorter100|14329_ ;
  assign \new_Sorter100|14429_  = \new_Sorter100|14328_  | \new_Sorter100|14329_ ;
  assign \new_Sorter100|14430_  = \new_Sorter100|14330_  & \new_Sorter100|14331_ ;
  assign \new_Sorter100|14431_  = \new_Sorter100|14330_  | \new_Sorter100|14331_ ;
  assign \new_Sorter100|14432_  = \new_Sorter100|14332_  & \new_Sorter100|14333_ ;
  assign \new_Sorter100|14433_  = \new_Sorter100|14332_  | \new_Sorter100|14333_ ;
  assign \new_Sorter100|14434_  = \new_Sorter100|14334_  & \new_Sorter100|14335_ ;
  assign \new_Sorter100|14435_  = \new_Sorter100|14334_  | \new_Sorter100|14335_ ;
  assign \new_Sorter100|14436_  = \new_Sorter100|14336_  & \new_Sorter100|14337_ ;
  assign \new_Sorter100|14437_  = \new_Sorter100|14336_  | \new_Sorter100|14337_ ;
  assign \new_Sorter100|14438_  = \new_Sorter100|14338_  & \new_Sorter100|14339_ ;
  assign \new_Sorter100|14439_  = \new_Sorter100|14338_  | \new_Sorter100|14339_ ;
  assign \new_Sorter100|14440_  = \new_Sorter100|14340_  & \new_Sorter100|14341_ ;
  assign \new_Sorter100|14441_  = \new_Sorter100|14340_  | \new_Sorter100|14341_ ;
  assign \new_Sorter100|14442_  = \new_Sorter100|14342_  & \new_Sorter100|14343_ ;
  assign \new_Sorter100|14443_  = \new_Sorter100|14342_  | \new_Sorter100|14343_ ;
  assign \new_Sorter100|14444_  = \new_Sorter100|14344_  & \new_Sorter100|14345_ ;
  assign \new_Sorter100|14445_  = \new_Sorter100|14344_  | \new_Sorter100|14345_ ;
  assign \new_Sorter100|14446_  = \new_Sorter100|14346_  & \new_Sorter100|14347_ ;
  assign \new_Sorter100|14447_  = \new_Sorter100|14346_  | \new_Sorter100|14347_ ;
  assign \new_Sorter100|14448_  = \new_Sorter100|14348_  & \new_Sorter100|14349_ ;
  assign \new_Sorter100|14449_  = \new_Sorter100|14348_  | \new_Sorter100|14349_ ;
  assign \new_Sorter100|14450_  = \new_Sorter100|14350_  & \new_Sorter100|14351_ ;
  assign \new_Sorter100|14451_  = \new_Sorter100|14350_  | \new_Sorter100|14351_ ;
  assign \new_Sorter100|14452_  = \new_Sorter100|14352_  & \new_Sorter100|14353_ ;
  assign \new_Sorter100|14453_  = \new_Sorter100|14352_  | \new_Sorter100|14353_ ;
  assign \new_Sorter100|14454_  = \new_Sorter100|14354_  & \new_Sorter100|14355_ ;
  assign \new_Sorter100|14455_  = \new_Sorter100|14354_  | \new_Sorter100|14355_ ;
  assign \new_Sorter100|14456_  = \new_Sorter100|14356_  & \new_Sorter100|14357_ ;
  assign \new_Sorter100|14457_  = \new_Sorter100|14356_  | \new_Sorter100|14357_ ;
  assign \new_Sorter100|14458_  = \new_Sorter100|14358_  & \new_Sorter100|14359_ ;
  assign \new_Sorter100|14459_  = \new_Sorter100|14358_  | \new_Sorter100|14359_ ;
  assign \new_Sorter100|14460_  = \new_Sorter100|14360_  & \new_Sorter100|14361_ ;
  assign \new_Sorter100|14461_  = \new_Sorter100|14360_  | \new_Sorter100|14361_ ;
  assign \new_Sorter100|14462_  = \new_Sorter100|14362_  & \new_Sorter100|14363_ ;
  assign \new_Sorter100|14463_  = \new_Sorter100|14362_  | \new_Sorter100|14363_ ;
  assign \new_Sorter100|14464_  = \new_Sorter100|14364_  & \new_Sorter100|14365_ ;
  assign \new_Sorter100|14465_  = \new_Sorter100|14364_  | \new_Sorter100|14365_ ;
  assign \new_Sorter100|14466_  = \new_Sorter100|14366_  & \new_Sorter100|14367_ ;
  assign \new_Sorter100|14467_  = \new_Sorter100|14366_  | \new_Sorter100|14367_ ;
  assign \new_Sorter100|14468_  = \new_Sorter100|14368_  & \new_Sorter100|14369_ ;
  assign \new_Sorter100|14469_  = \new_Sorter100|14368_  | \new_Sorter100|14369_ ;
  assign \new_Sorter100|14470_  = \new_Sorter100|14370_  & \new_Sorter100|14371_ ;
  assign \new_Sorter100|14471_  = \new_Sorter100|14370_  | \new_Sorter100|14371_ ;
  assign \new_Sorter100|14472_  = \new_Sorter100|14372_  & \new_Sorter100|14373_ ;
  assign \new_Sorter100|14473_  = \new_Sorter100|14372_  | \new_Sorter100|14373_ ;
  assign \new_Sorter100|14474_  = \new_Sorter100|14374_  & \new_Sorter100|14375_ ;
  assign \new_Sorter100|14475_  = \new_Sorter100|14374_  | \new_Sorter100|14375_ ;
  assign \new_Sorter100|14476_  = \new_Sorter100|14376_  & \new_Sorter100|14377_ ;
  assign \new_Sorter100|14477_  = \new_Sorter100|14376_  | \new_Sorter100|14377_ ;
  assign \new_Sorter100|14478_  = \new_Sorter100|14378_  & \new_Sorter100|14379_ ;
  assign \new_Sorter100|14479_  = \new_Sorter100|14378_  | \new_Sorter100|14379_ ;
  assign \new_Sorter100|14480_  = \new_Sorter100|14380_  & \new_Sorter100|14381_ ;
  assign \new_Sorter100|14481_  = \new_Sorter100|14380_  | \new_Sorter100|14381_ ;
  assign \new_Sorter100|14482_  = \new_Sorter100|14382_  & \new_Sorter100|14383_ ;
  assign \new_Sorter100|14483_  = \new_Sorter100|14382_  | \new_Sorter100|14383_ ;
  assign \new_Sorter100|14484_  = \new_Sorter100|14384_  & \new_Sorter100|14385_ ;
  assign \new_Sorter100|14485_  = \new_Sorter100|14384_  | \new_Sorter100|14385_ ;
  assign \new_Sorter100|14486_  = \new_Sorter100|14386_  & \new_Sorter100|14387_ ;
  assign \new_Sorter100|14487_  = \new_Sorter100|14386_  | \new_Sorter100|14387_ ;
  assign \new_Sorter100|14488_  = \new_Sorter100|14388_  & \new_Sorter100|14389_ ;
  assign \new_Sorter100|14489_  = \new_Sorter100|14388_  | \new_Sorter100|14389_ ;
  assign \new_Sorter100|14490_  = \new_Sorter100|14390_  & \new_Sorter100|14391_ ;
  assign \new_Sorter100|14491_  = \new_Sorter100|14390_  | \new_Sorter100|14391_ ;
  assign \new_Sorter100|14492_  = \new_Sorter100|14392_  & \new_Sorter100|14393_ ;
  assign \new_Sorter100|14493_  = \new_Sorter100|14392_  | \new_Sorter100|14393_ ;
  assign \new_Sorter100|14494_  = \new_Sorter100|14394_  & \new_Sorter100|14395_ ;
  assign \new_Sorter100|14495_  = \new_Sorter100|14394_  | \new_Sorter100|14395_ ;
  assign \new_Sorter100|14496_  = \new_Sorter100|14396_  & \new_Sorter100|14397_ ;
  assign \new_Sorter100|14497_  = \new_Sorter100|14396_  | \new_Sorter100|14397_ ;
  assign \new_Sorter100|14498_  = \new_Sorter100|14398_  & \new_Sorter100|14399_ ;
  assign \new_Sorter100|14499_  = \new_Sorter100|14398_  | \new_Sorter100|14399_ ;
  assign \new_Sorter100|14500_  = \new_Sorter100|14400_ ;
  assign \new_Sorter100|14599_  = \new_Sorter100|14499_ ;
  assign \new_Sorter100|14501_  = \new_Sorter100|14401_  & \new_Sorter100|14402_ ;
  assign \new_Sorter100|14502_  = \new_Sorter100|14401_  | \new_Sorter100|14402_ ;
  assign \new_Sorter100|14503_  = \new_Sorter100|14403_  & \new_Sorter100|14404_ ;
  assign \new_Sorter100|14504_  = \new_Sorter100|14403_  | \new_Sorter100|14404_ ;
  assign \new_Sorter100|14505_  = \new_Sorter100|14405_  & \new_Sorter100|14406_ ;
  assign \new_Sorter100|14506_  = \new_Sorter100|14405_  | \new_Sorter100|14406_ ;
  assign \new_Sorter100|14507_  = \new_Sorter100|14407_  & \new_Sorter100|14408_ ;
  assign \new_Sorter100|14508_  = \new_Sorter100|14407_  | \new_Sorter100|14408_ ;
  assign \new_Sorter100|14509_  = \new_Sorter100|14409_  & \new_Sorter100|14410_ ;
  assign \new_Sorter100|14510_  = \new_Sorter100|14409_  | \new_Sorter100|14410_ ;
  assign \new_Sorter100|14511_  = \new_Sorter100|14411_  & \new_Sorter100|14412_ ;
  assign \new_Sorter100|14512_  = \new_Sorter100|14411_  | \new_Sorter100|14412_ ;
  assign \new_Sorter100|14513_  = \new_Sorter100|14413_  & \new_Sorter100|14414_ ;
  assign \new_Sorter100|14514_  = \new_Sorter100|14413_  | \new_Sorter100|14414_ ;
  assign \new_Sorter100|14515_  = \new_Sorter100|14415_  & \new_Sorter100|14416_ ;
  assign \new_Sorter100|14516_  = \new_Sorter100|14415_  | \new_Sorter100|14416_ ;
  assign \new_Sorter100|14517_  = \new_Sorter100|14417_  & \new_Sorter100|14418_ ;
  assign \new_Sorter100|14518_  = \new_Sorter100|14417_  | \new_Sorter100|14418_ ;
  assign \new_Sorter100|14519_  = \new_Sorter100|14419_  & \new_Sorter100|14420_ ;
  assign \new_Sorter100|14520_  = \new_Sorter100|14419_  | \new_Sorter100|14420_ ;
  assign \new_Sorter100|14521_  = \new_Sorter100|14421_  & \new_Sorter100|14422_ ;
  assign \new_Sorter100|14522_  = \new_Sorter100|14421_  | \new_Sorter100|14422_ ;
  assign \new_Sorter100|14523_  = \new_Sorter100|14423_  & \new_Sorter100|14424_ ;
  assign \new_Sorter100|14524_  = \new_Sorter100|14423_  | \new_Sorter100|14424_ ;
  assign \new_Sorter100|14525_  = \new_Sorter100|14425_  & \new_Sorter100|14426_ ;
  assign \new_Sorter100|14526_  = \new_Sorter100|14425_  | \new_Sorter100|14426_ ;
  assign \new_Sorter100|14527_  = \new_Sorter100|14427_  & \new_Sorter100|14428_ ;
  assign \new_Sorter100|14528_  = \new_Sorter100|14427_  | \new_Sorter100|14428_ ;
  assign \new_Sorter100|14529_  = \new_Sorter100|14429_  & \new_Sorter100|14430_ ;
  assign \new_Sorter100|14530_  = \new_Sorter100|14429_  | \new_Sorter100|14430_ ;
  assign \new_Sorter100|14531_  = \new_Sorter100|14431_  & \new_Sorter100|14432_ ;
  assign \new_Sorter100|14532_  = \new_Sorter100|14431_  | \new_Sorter100|14432_ ;
  assign \new_Sorter100|14533_  = \new_Sorter100|14433_  & \new_Sorter100|14434_ ;
  assign \new_Sorter100|14534_  = \new_Sorter100|14433_  | \new_Sorter100|14434_ ;
  assign \new_Sorter100|14535_  = \new_Sorter100|14435_  & \new_Sorter100|14436_ ;
  assign \new_Sorter100|14536_  = \new_Sorter100|14435_  | \new_Sorter100|14436_ ;
  assign \new_Sorter100|14537_  = \new_Sorter100|14437_  & \new_Sorter100|14438_ ;
  assign \new_Sorter100|14538_  = \new_Sorter100|14437_  | \new_Sorter100|14438_ ;
  assign \new_Sorter100|14539_  = \new_Sorter100|14439_  & \new_Sorter100|14440_ ;
  assign \new_Sorter100|14540_  = \new_Sorter100|14439_  | \new_Sorter100|14440_ ;
  assign \new_Sorter100|14541_  = \new_Sorter100|14441_  & \new_Sorter100|14442_ ;
  assign \new_Sorter100|14542_  = \new_Sorter100|14441_  | \new_Sorter100|14442_ ;
  assign \new_Sorter100|14543_  = \new_Sorter100|14443_  & \new_Sorter100|14444_ ;
  assign \new_Sorter100|14544_  = \new_Sorter100|14443_  | \new_Sorter100|14444_ ;
  assign \new_Sorter100|14545_  = \new_Sorter100|14445_  & \new_Sorter100|14446_ ;
  assign \new_Sorter100|14546_  = \new_Sorter100|14445_  | \new_Sorter100|14446_ ;
  assign \new_Sorter100|14547_  = \new_Sorter100|14447_  & \new_Sorter100|14448_ ;
  assign \new_Sorter100|14548_  = \new_Sorter100|14447_  | \new_Sorter100|14448_ ;
  assign \new_Sorter100|14549_  = \new_Sorter100|14449_  & \new_Sorter100|14450_ ;
  assign \new_Sorter100|14550_  = \new_Sorter100|14449_  | \new_Sorter100|14450_ ;
  assign \new_Sorter100|14551_  = \new_Sorter100|14451_  & \new_Sorter100|14452_ ;
  assign \new_Sorter100|14552_  = \new_Sorter100|14451_  | \new_Sorter100|14452_ ;
  assign \new_Sorter100|14553_  = \new_Sorter100|14453_  & \new_Sorter100|14454_ ;
  assign \new_Sorter100|14554_  = \new_Sorter100|14453_  | \new_Sorter100|14454_ ;
  assign \new_Sorter100|14555_  = \new_Sorter100|14455_  & \new_Sorter100|14456_ ;
  assign \new_Sorter100|14556_  = \new_Sorter100|14455_  | \new_Sorter100|14456_ ;
  assign \new_Sorter100|14557_  = \new_Sorter100|14457_  & \new_Sorter100|14458_ ;
  assign \new_Sorter100|14558_  = \new_Sorter100|14457_  | \new_Sorter100|14458_ ;
  assign \new_Sorter100|14559_  = \new_Sorter100|14459_  & \new_Sorter100|14460_ ;
  assign \new_Sorter100|14560_  = \new_Sorter100|14459_  | \new_Sorter100|14460_ ;
  assign \new_Sorter100|14561_  = \new_Sorter100|14461_  & \new_Sorter100|14462_ ;
  assign \new_Sorter100|14562_  = \new_Sorter100|14461_  | \new_Sorter100|14462_ ;
  assign \new_Sorter100|14563_  = \new_Sorter100|14463_  & \new_Sorter100|14464_ ;
  assign \new_Sorter100|14564_  = \new_Sorter100|14463_  | \new_Sorter100|14464_ ;
  assign \new_Sorter100|14565_  = \new_Sorter100|14465_  & \new_Sorter100|14466_ ;
  assign \new_Sorter100|14566_  = \new_Sorter100|14465_  | \new_Sorter100|14466_ ;
  assign \new_Sorter100|14567_  = \new_Sorter100|14467_  & \new_Sorter100|14468_ ;
  assign \new_Sorter100|14568_  = \new_Sorter100|14467_  | \new_Sorter100|14468_ ;
  assign \new_Sorter100|14569_  = \new_Sorter100|14469_  & \new_Sorter100|14470_ ;
  assign \new_Sorter100|14570_  = \new_Sorter100|14469_  | \new_Sorter100|14470_ ;
  assign \new_Sorter100|14571_  = \new_Sorter100|14471_  & \new_Sorter100|14472_ ;
  assign \new_Sorter100|14572_  = \new_Sorter100|14471_  | \new_Sorter100|14472_ ;
  assign \new_Sorter100|14573_  = \new_Sorter100|14473_  & \new_Sorter100|14474_ ;
  assign \new_Sorter100|14574_  = \new_Sorter100|14473_  | \new_Sorter100|14474_ ;
  assign \new_Sorter100|14575_  = \new_Sorter100|14475_  & \new_Sorter100|14476_ ;
  assign \new_Sorter100|14576_  = \new_Sorter100|14475_  | \new_Sorter100|14476_ ;
  assign \new_Sorter100|14577_  = \new_Sorter100|14477_  & \new_Sorter100|14478_ ;
  assign \new_Sorter100|14578_  = \new_Sorter100|14477_  | \new_Sorter100|14478_ ;
  assign \new_Sorter100|14579_  = \new_Sorter100|14479_  & \new_Sorter100|14480_ ;
  assign \new_Sorter100|14580_  = \new_Sorter100|14479_  | \new_Sorter100|14480_ ;
  assign \new_Sorter100|14581_  = \new_Sorter100|14481_  & \new_Sorter100|14482_ ;
  assign \new_Sorter100|14582_  = \new_Sorter100|14481_  | \new_Sorter100|14482_ ;
  assign \new_Sorter100|14583_  = \new_Sorter100|14483_  & \new_Sorter100|14484_ ;
  assign \new_Sorter100|14584_  = \new_Sorter100|14483_  | \new_Sorter100|14484_ ;
  assign \new_Sorter100|14585_  = \new_Sorter100|14485_  & \new_Sorter100|14486_ ;
  assign \new_Sorter100|14586_  = \new_Sorter100|14485_  | \new_Sorter100|14486_ ;
  assign \new_Sorter100|14587_  = \new_Sorter100|14487_  & \new_Sorter100|14488_ ;
  assign \new_Sorter100|14588_  = \new_Sorter100|14487_  | \new_Sorter100|14488_ ;
  assign \new_Sorter100|14589_  = \new_Sorter100|14489_  & \new_Sorter100|14490_ ;
  assign \new_Sorter100|14590_  = \new_Sorter100|14489_  | \new_Sorter100|14490_ ;
  assign \new_Sorter100|14591_  = \new_Sorter100|14491_  & \new_Sorter100|14492_ ;
  assign \new_Sorter100|14592_  = \new_Sorter100|14491_  | \new_Sorter100|14492_ ;
  assign \new_Sorter100|14593_  = \new_Sorter100|14493_  & \new_Sorter100|14494_ ;
  assign \new_Sorter100|14594_  = \new_Sorter100|14493_  | \new_Sorter100|14494_ ;
  assign \new_Sorter100|14595_  = \new_Sorter100|14495_  & \new_Sorter100|14496_ ;
  assign \new_Sorter100|14596_  = \new_Sorter100|14495_  | \new_Sorter100|14496_ ;
  assign \new_Sorter100|14597_  = \new_Sorter100|14497_  & \new_Sorter100|14498_ ;
  assign \new_Sorter100|14598_  = \new_Sorter100|14497_  | \new_Sorter100|14498_ ;
  assign \new_Sorter100|14600_  = \new_Sorter100|14500_  & \new_Sorter100|14501_ ;
  assign \new_Sorter100|14601_  = \new_Sorter100|14500_  | \new_Sorter100|14501_ ;
  assign \new_Sorter100|14602_  = \new_Sorter100|14502_  & \new_Sorter100|14503_ ;
  assign \new_Sorter100|14603_  = \new_Sorter100|14502_  | \new_Sorter100|14503_ ;
  assign \new_Sorter100|14604_  = \new_Sorter100|14504_  & \new_Sorter100|14505_ ;
  assign \new_Sorter100|14605_  = \new_Sorter100|14504_  | \new_Sorter100|14505_ ;
  assign \new_Sorter100|14606_  = \new_Sorter100|14506_  & \new_Sorter100|14507_ ;
  assign \new_Sorter100|14607_  = \new_Sorter100|14506_  | \new_Sorter100|14507_ ;
  assign \new_Sorter100|14608_  = \new_Sorter100|14508_  & \new_Sorter100|14509_ ;
  assign \new_Sorter100|14609_  = \new_Sorter100|14508_  | \new_Sorter100|14509_ ;
  assign \new_Sorter100|14610_  = \new_Sorter100|14510_  & \new_Sorter100|14511_ ;
  assign \new_Sorter100|14611_  = \new_Sorter100|14510_  | \new_Sorter100|14511_ ;
  assign \new_Sorter100|14612_  = \new_Sorter100|14512_  & \new_Sorter100|14513_ ;
  assign \new_Sorter100|14613_  = \new_Sorter100|14512_  | \new_Sorter100|14513_ ;
  assign \new_Sorter100|14614_  = \new_Sorter100|14514_  & \new_Sorter100|14515_ ;
  assign \new_Sorter100|14615_  = \new_Sorter100|14514_  | \new_Sorter100|14515_ ;
  assign \new_Sorter100|14616_  = \new_Sorter100|14516_  & \new_Sorter100|14517_ ;
  assign \new_Sorter100|14617_  = \new_Sorter100|14516_  | \new_Sorter100|14517_ ;
  assign \new_Sorter100|14618_  = \new_Sorter100|14518_  & \new_Sorter100|14519_ ;
  assign \new_Sorter100|14619_  = \new_Sorter100|14518_  | \new_Sorter100|14519_ ;
  assign \new_Sorter100|14620_  = \new_Sorter100|14520_  & \new_Sorter100|14521_ ;
  assign \new_Sorter100|14621_  = \new_Sorter100|14520_  | \new_Sorter100|14521_ ;
  assign \new_Sorter100|14622_  = \new_Sorter100|14522_  & \new_Sorter100|14523_ ;
  assign \new_Sorter100|14623_  = \new_Sorter100|14522_  | \new_Sorter100|14523_ ;
  assign \new_Sorter100|14624_  = \new_Sorter100|14524_  & \new_Sorter100|14525_ ;
  assign \new_Sorter100|14625_  = \new_Sorter100|14524_  | \new_Sorter100|14525_ ;
  assign \new_Sorter100|14626_  = \new_Sorter100|14526_  & \new_Sorter100|14527_ ;
  assign \new_Sorter100|14627_  = \new_Sorter100|14526_  | \new_Sorter100|14527_ ;
  assign \new_Sorter100|14628_  = \new_Sorter100|14528_  & \new_Sorter100|14529_ ;
  assign \new_Sorter100|14629_  = \new_Sorter100|14528_  | \new_Sorter100|14529_ ;
  assign \new_Sorter100|14630_  = \new_Sorter100|14530_  & \new_Sorter100|14531_ ;
  assign \new_Sorter100|14631_  = \new_Sorter100|14530_  | \new_Sorter100|14531_ ;
  assign \new_Sorter100|14632_  = \new_Sorter100|14532_  & \new_Sorter100|14533_ ;
  assign \new_Sorter100|14633_  = \new_Sorter100|14532_  | \new_Sorter100|14533_ ;
  assign \new_Sorter100|14634_  = \new_Sorter100|14534_  & \new_Sorter100|14535_ ;
  assign \new_Sorter100|14635_  = \new_Sorter100|14534_  | \new_Sorter100|14535_ ;
  assign \new_Sorter100|14636_  = \new_Sorter100|14536_  & \new_Sorter100|14537_ ;
  assign \new_Sorter100|14637_  = \new_Sorter100|14536_  | \new_Sorter100|14537_ ;
  assign \new_Sorter100|14638_  = \new_Sorter100|14538_  & \new_Sorter100|14539_ ;
  assign \new_Sorter100|14639_  = \new_Sorter100|14538_  | \new_Sorter100|14539_ ;
  assign \new_Sorter100|14640_  = \new_Sorter100|14540_  & \new_Sorter100|14541_ ;
  assign \new_Sorter100|14641_  = \new_Sorter100|14540_  | \new_Sorter100|14541_ ;
  assign \new_Sorter100|14642_  = \new_Sorter100|14542_  & \new_Sorter100|14543_ ;
  assign \new_Sorter100|14643_  = \new_Sorter100|14542_  | \new_Sorter100|14543_ ;
  assign \new_Sorter100|14644_  = \new_Sorter100|14544_  & \new_Sorter100|14545_ ;
  assign \new_Sorter100|14645_  = \new_Sorter100|14544_  | \new_Sorter100|14545_ ;
  assign \new_Sorter100|14646_  = \new_Sorter100|14546_  & \new_Sorter100|14547_ ;
  assign \new_Sorter100|14647_  = \new_Sorter100|14546_  | \new_Sorter100|14547_ ;
  assign \new_Sorter100|14648_  = \new_Sorter100|14548_  & \new_Sorter100|14549_ ;
  assign \new_Sorter100|14649_  = \new_Sorter100|14548_  | \new_Sorter100|14549_ ;
  assign \new_Sorter100|14650_  = \new_Sorter100|14550_  & \new_Sorter100|14551_ ;
  assign \new_Sorter100|14651_  = \new_Sorter100|14550_  | \new_Sorter100|14551_ ;
  assign \new_Sorter100|14652_  = \new_Sorter100|14552_  & \new_Sorter100|14553_ ;
  assign \new_Sorter100|14653_  = \new_Sorter100|14552_  | \new_Sorter100|14553_ ;
  assign \new_Sorter100|14654_  = \new_Sorter100|14554_  & \new_Sorter100|14555_ ;
  assign \new_Sorter100|14655_  = \new_Sorter100|14554_  | \new_Sorter100|14555_ ;
  assign \new_Sorter100|14656_  = \new_Sorter100|14556_  & \new_Sorter100|14557_ ;
  assign \new_Sorter100|14657_  = \new_Sorter100|14556_  | \new_Sorter100|14557_ ;
  assign \new_Sorter100|14658_  = \new_Sorter100|14558_  & \new_Sorter100|14559_ ;
  assign \new_Sorter100|14659_  = \new_Sorter100|14558_  | \new_Sorter100|14559_ ;
  assign \new_Sorter100|14660_  = \new_Sorter100|14560_  & \new_Sorter100|14561_ ;
  assign \new_Sorter100|14661_  = \new_Sorter100|14560_  | \new_Sorter100|14561_ ;
  assign \new_Sorter100|14662_  = \new_Sorter100|14562_  & \new_Sorter100|14563_ ;
  assign \new_Sorter100|14663_  = \new_Sorter100|14562_  | \new_Sorter100|14563_ ;
  assign \new_Sorter100|14664_  = \new_Sorter100|14564_  & \new_Sorter100|14565_ ;
  assign \new_Sorter100|14665_  = \new_Sorter100|14564_  | \new_Sorter100|14565_ ;
  assign \new_Sorter100|14666_  = \new_Sorter100|14566_  & \new_Sorter100|14567_ ;
  assign \new_Sorter100|14667_  = \new_Sorter100|14566_  | \new_Sorter100|14567_ ;
  assign \new_Sorter100|14668_  = \new_Sorter100|14568_  & \new_Sorter100|14569_ ;
  assign \new_Sorter100|14669_  = \new_Sorter100|14568_  | \new_Sorter100|14569_ ;
  assign \new_Sorter100|14670_  = \new_Sorter100|14570_  & \new_Sorter100|14571_ ;
  assign \new_Sorter100|14671_  = \new_Sorter100|14570_  | \new_Sorter100|14571_ ;
  assign \new_Sorter100|14672_  = \new_Sorter100|14572_  & \new_Sorter100|14573_ ;
  assign \new_Sorter100|14673_  = \new_Sorter100|14572_  | \new_Sorter100|14573_ ;
  assign \new_Sorter100|14674_  = \new_Sorter100|14574_  & \new_Sorter100|14575_ ;
  assign \new_Sorter100|14675_  = \new_Sorter100|14574_  | \new_Sorter100|14575_ ;
  assign \new_Sorter100|14676_  = \new_Sorter100|14576_  & \new_Sorter100|14577_ ;
  assign \new_Sorter100|14677_  = \new_Sorter100|14576_  | \new_Sorter100|14577_ ;
  assign \new_Sorter100|14678_  = \new_Sorter100|14578_  & \new_Sorter100|14579_ ;
  assign \new_Sorter100|14679_  = \new_Sorter100|14578_  | \new_Sorter100|14579_ ;
  assign \new_Sorter100|14680_  = \new_Sorter100|14580_  & \new_Sorter100|14581_ ;
  assign \new_Sorter100|14681_  = \new_Sorter100|14580_  | \new_Sorter100|14581_ ;
  assign \new_Sorter100|14682_  = \new_Sorter100|14582_  & \new_Sorter100|14583_ ;
  assign \new_Sorter100|14683_  = \new_Sorter100|14582_  | \new_Sorter100|14583_ ;
  assign \new_Sorter100|14684_  = \new_Sorter100|14584_  & \new_Sorter100|14585_ ;
  assign \new_Sorter100|14685_  = \new_Sorter100|14584_  | \new_Sorter100|14585_ ;
  assign \new_Sorter100|14686_  = \new_Sorter100|14586_  & \new_Sorter100|14587_ ;
  assign \new_Sorter100|14687_  = \new_Sorter100|14586_  | \new_Sorter100|14587_ ;
  assign \new_Sorter100|14688_  = \new_Sorter100|14588_  & \new_Sorter100|14589_ ;
  assign \new_Sorter100|14689_  = \new_Sorter100|14588_  | \new_Sorter100|14589_ ;
  assign \new_Sorter100|14690_  = \new_Sorter100|14590_  & \new_Sorter100|14591_ ;
  assign \new_Sorter100|14691_  = \new_Sorter100|14590_  | \new_Sorter100|14591_ ;
  assign \new_Sorter100|14692_  = \new_Sorter100|14592_  & \new_Sorter100|14593_ ;
  assign \new_Sorter100|14693_  = \new_Sorter100|14592_  | \new_Sorter100|14593_ ;
  assign \new_Sorter100|14694_  = \new_Sorter100|14594_  & \new_Sorter100|14595_ ;
  assign \new_Sorter100|14695_  = \new_Sorter100|14594_  | \new_Sorter100|14595_ ;
  assign \new_Sorter100|14696_  = \new_Sorter100|14596_  & \new_Sorter100|14597_ ;
  assign \new_Sorter100|14697_  = \new_Sorter100|14596_  | \new_Sorter100|14597_ ;
  assign \new_Sorter100|14698_  = \new_Sorter100|14598_  & \new_Sorter100|14599_ ;
  assign \new_Sorter100|14699_  = \new_Sorter100|14598_  | \new_Sorter100|14599_ ;
  assign \new_Sorter100|14700_  = \new_Sorter100|14600_ ;
  assign \new_Sorter100|14799_  = \new_Sorter100|14699_ ;
  assign \new_Sorter100|14701_  = \new_Sorter100|14601_  & \new_Sorter100|14602_ ;
  assign \new_Sorter100|14702_  = \new_Sorter100|14601_  | \new_Sorter100|14602_ ;
  assign \new_Sorter100|14703_  = \new_Sorter100|14603_  & \new_Sorter100|14604_ ;
  assign \new_Sorter100|14704_  = \new_Sorter100|14603_  | \new_Sorter100|14604_ ;
  assign \new_Sorter100|14705_  = \new_Sorter100|14605_  & \new_Sorter100|14606_ ;
  assign \new_Sorter100|14706_  = \new_Sorter100|14605_  | \new_Sorter100|14606_ ;
  assign \new_Sorter100|14707_  = \new_Sorter100|14607_  & \new_Sorter100|14608_ ;
  assign \new_Sorter100|14708_  = \new_Sorter100|14607_  | \new_Sorter100|14608_ ;
  assign \new_Sorter100|14709_  = \new_Sorter100|14609_  & \new_Sorter100|14610_ ;
  assign \new_Sorter100|14710_  = \new_Sorter100|14609_  | \new_Sorter100|14610_ ;
  assign \new_Sorter100|14711_  = \new_Sorter100|14611_  & \new_Sorter100|14612_ ;
  assign \new_Sorter100|14712_  = \new_Sorter100|14611_  | \new_Sorter100|14612_ ;
  assign \new_Sorter100|14713_  = \new_Sorter100|14613_  & \new_Sorter100|14614_ ;
  assign \new_Sorter100|14714_  = \new_Sorter100|14613_  | \new_Sorter100|14614_ ;
  assign \new_Sorter100|14715_  = \new_Sorter100|14615_  & \new_Sorter100|14616_ ;
  assign \new_Sorter100|14716_  = \new_Sorter100|14615_  | \new_Sorter100|14616_ ;
  assign \new_Sorter100|14717_  = \new_Sorter100|14617_  & \new_Sorter100|14618_ ;
  assign \new_Sorter100|14718_  = \new_Sorter100|14617_  | \new_Sorter100|14618_ ;
  assign \new_Sorter100|14719_  = \new_Sorter100|14619_  & \new_Sorter100|14620_ ;
  assign \new_Sorter100|14720_  = \new_Sorter100|14619_  | \new_Sorter100|14620_ ;
  assign \new_Sorter100|14721_  = \new_Sorter100|14621_  & \new_Sorter100|14622_ ;
  assign \new_Sorter100|14722_  = \new_Sorter100|14621_  | \new_Sorter100|14622_ ;
  assign \new_Sorter100|14723_  = \new_Sorter100|14623_  & \new_Sorter100|14624_ ;
  assign \new_Sorter100|14724_  = \new_Sorter100|14623_  | \new_Sorter100|14624_ ;
  assign \new_Sorter100|14725_  = \new_Sorter100|14625_  & \new_Sorter100|14626_ ;
  assign \new_Sorter100|14726_  = \new_Sorter100|14625_  | \new_Sorter100|14626_ ;
  assign \new_Sorter100|14727_  = \new_Sorter100|14627_  & \new_Sorter100|14628_ ;
  assign \new_Sorter100|14728_  = \new_Sorter100|14627_  | \new_Sorter100|14628_ ;
  assign \new_Sorter100|14729_  = \new_Sorter100|14629_  & \new_Sorter100|14630_ ;
  assign \new_Sorter100|14730_  = \new_Sorter100|14629_  | \new_Sorter100|14630_ ;
  assign \new_Sorter100|14731_  = \new_Sorter100|14631_  & \new_Sorter100|14632_ ;
  assign \new_Sorter100|14732_  = \new_Sorter100|14631_  | \new_Sorter100|14632_ ;
  assign \new_Sorter100|14733_  = \new_Sorter100|14633_  & \new_Sorter100|14634_ ;
  assign \new_Sorter100|14734_  = \new_Sorter100|14633_  | \new_Sorter100|14634_ ;
  assign \new_Sorter100|14735_  = \new_Sorter100|14635_  & \new_Sorter100|14636_ ;
  assign \new_Sorter100|14736_  = \new_Sorter100|14635_  | \new_Sorter100|14636_ ;
  assign \new_Sorter100|14737_  = \new_Sorter100|14637_  & \new_Sorter100|14638_ ;
  assign \new_Sorter100|14738_  = \new_Sorter100|14637_  | \new_Sorter100|14638_ ;
  assign \new_Sorter100|14739_  = \new_Sorter100|14639_  & \new_Sorter100|14640_ ;
  assign \new_Sorter100|14740_  = \new_Sorter100|14639_  | \new_Sorter100|14640_ ;
  assign \new_Sorter100|14741_  = \new_Sorter100|14641_  & \new_Sorter100|14642_ ;
  assign \new_Sorter100|14742_  = \new_Sorter100|14641_  | \new_Sorter100|14642_ ;
  assign \new_Sorter100|14743_  = \new_Sorter100|14643_  & \new_Sorter100|14644_ ;
  assign \new_Sorter100|14744_  = \new_Sorter100|14643_  | \new_Sorter100|14644_ ;
  assign \new_Sorter100|14745_  = \new_Sorter100|14645_  & \new_Sorter100|14646_ ;
  assign \new_Sorter100|14746_  = \new_Sorter100|14645_  | \new_Sorter100|14646_ ;
  assign \new_Sorter100|14747_  = \new_Sorter100|14647_  & \new_Sorter100|14648_ ;
  assign \new_Sorter100|14748_  = \new_Sorter100|14647_  | \new_Sorter100|14648_ ;
  assign \new_Sorter100|14749_  = \new_Sorter100|14649_  & \new_Sorter100|14650_ ;
  assign \new_Sorter100|14750_  = \new_Sorter100|14649_  | \new_Sorter100|14650_ ;
  assign \new_Sorter100|14751_  = \new_Sorter100|14651_  & \new_Sorter100|14652_ ;
  assign \new_Sorter100|14752_  = \new_Sorter100|14651_  | \new_Sorter100|14652_ ;
  assign \new_Sorter100|14753_  = \new_Sorter100|14653_  & \new_Sorter100|14654_ ;
  assign \new_Sorter100|14754_  = \new_Sorter100|14653_  | \new_Sorter100|14654_ ;
  assign \new_Sorter100|14755_  = \new_Sorter100|14655_  & \new_Sorter100|14656_ ;
  assign \new_Sorter100|14756_  = \new_Sorter100|14655_  | \new_Sorter100|14656_ ;
  assign \new_Sorter100|14757_  = \new_Sorter100|14657_  & \new_Sorter100|14658_ ;
  assign \new_Sorter100|14758_  = \new_Sorter100|14657_  | \new_Sorter100|14658_ ;
  assign \new_Sorter100|14759_  = \new_Sorter100|14659_  & \new_Sorter100|14660_ ;
  assign \new_Sorter100|14760_  = \new_Sorter100|14659_  | \new_Sorter100|14660_ ;
  assign \new_Sorter100|14761_  = \new_Sorter100|14661_  & \new_Sorter100|14662_ ;
  assign \new_Sorter100|14762_  = \new_Sorter100|14661_  | \new_Sorter100|14662_ ;
  assign \new_Sorter100|14763_  = \new_Sorter100|14663_  & \new_Sorter100|14664_ ;
  assign \new_Sorter100|14764_  = \new_Sorter100|14663_  | \new_Sorter100|14664_ ;
  assign \new_Sorter100|14765_  = \new_Sorter100|14665_  & \new_Sorter100|14666_ ;
  assign \new_Sorter100|14766_  = \new_Sorter100|14665_  | \new_Sorter100|14666_ ;
  assign \new_Sorter100|14767_  = \new_Sorter100|14667_  & \new_Sorter100|14668_ ;
  assign \new_Sorter100|14768_  = \new_Sorter100|14667_  | \new_Sorter100|14668_ ;
  assign \new_Sorter100|14769_  = \new_Sorter100|14669_  & \new_Sorter100|14670_ ;
  assign \new_Sorter100|14770_  = \new_Sorter100|14669_  | \new_Sorter100|14670_ ;
  assign \new_Sorter100|14771_  = \new_Sorter100|14671_  & \new_Sorter100|14672_ ;
  assign \new_Sorter100|14772_  = \new_Sorter100|14671_  | \new_Sorter100|14672_ ;
  assign \new_Sorter100|14773_  = \new_Sorter100|14673_  & \new_Sorter100|14674_ ;
  assign \new_Sorter100|14774_  = \new_Sorter100|14673_  | \new_Sorter100|14674_ ;
  assign \new_Sorter100|14775_  = \new_Sorter100|14675_  & \new_Sorter100|14676_ ;
  assign \new_Sorter100|14776_  = \new_Sorter100|14675_  | \new_Sorter100|14676_ ;
  assign \new_Sorter100|14777_  = \new_Sorter100|14677_  & \new_Sorter100|14678_ ;
  assign \new_Sorter100|14778_  = \new_Sorter100|14677_  | \new_Sorter100|14678_ ;
  assign \new_Sorter100|14779_  = \new_Sorter100|14679_  & \new_Sorter100|14680_ ;
  assign \new_Sorter100|14780_  = \new_Sorter100|14679_  | \new_Sorter100|14680_ ;
  assign \new_Sorter100|14781_  = \new_Sorter100|14681_  & \new_Sorter100|14682_ ;
  assign \new_Sorter100|14782_  = \new_Sorter100|14681_  | \new_Sorter100|14682_ ;
  assign \new_Sorter100|14783_  = \new_Sorter100|14683_  & \new_Sorter100|14684_ ;
  assign \new_Sorter100|14784_  = \new_Sorter100|14683_  | \new_Sorter100|14684_ ;
  assign \new_Sorter100|14785_  = \new_Sorter100|14685_  & \new_Sorter100|14686_ ;
  assign \new_Sorter100|14786_  = \new_Sorter100|14685_  | \new_Sorter100|14686_ ;
  assign \new_Sorter100|14787_  = \new_Sorter100|14687_  & \new_Sorter100|14688_ ;
  assign \new_Sorter100|14788_  = \new_Sorter100|14687_  | \new_Sorter100|14688_ ;
  assign \new_Sorter100|14789_  = \new_Sorter100|14689_  & \new_Sorter100|14690_ ;
  assign \new_Sorter100|14790_  = \new_Sorter100|14689_  | \new_Sorter100|14690_ ;
  assign \new_Sorter100|14791_  = \new_Sorter100|14691_  & \new_Sorter100|14692_ ;
  assign \new_Sorter100|14792_  = \new_Sorter100|14691_  | \new_Sorter100|14692_ ;
  assign \new_Sorter100|14793_  = \new_Sorter100|14693_  & \new_Sorter100|14694_ ;
  assign \new_Sorter100|14794_  = \new_Sorter100|14693_  | \new_Sorter100|14694_ ;
  assign \new_Sorter100|14795_  = \new_Sorter100|14695_  & \new_Sorter100|14696_ ;
  assign \new_Sorter100|14796_  = \new_Sorter100|14695_  | \new_Sorter100|14696_ ;
  assign \new_Sorter100|14797_  = \new_Sorter100|14697_  & \new_Sorter100|14698_ ;
  assign \new_Sorter100|14798_  = \new_Sorter100|14697_  | \new_Sorter100|14698_ ;
  assign \new_Sorter100|14800_  = \new_Sorter100|14700_  & \new_Sorter100|14701_ ;
  assign \new_Sorter100|14801_  = \new_Sorter100|14700_  | \new_Sorter100|14701_ ;
  assign \new_Sorter100|14802_  = \new_Sorter100|14702_  & \new_Sorter100|14703_ ;
  assign \new_Sorter100|14803_  = \new_Sorter100|14702_  | \new_Sorter100|14703_ ;
  assign \new_Sorter100|14804_  = \new_Sorter100|14704_  & \new_Sorter100|14705_ ;
  assign \new_Sorter100|14805_  = \new_Sorter100|14704_  | \new_Sorter100|14705_ ;
  assign \new_Sorter100|14806_  = \new_Sorter100|14706_  & \new_Sorter100|14707_ ;
  assign \new_Sorter100|14807_  = \new_Sorter100|14706_  | \new_Sorter100|14707_ ;
  assign \new_Sorter100|14808_  = \new_Sorter100|14708_  & \new_Sorter100|14709_ ;
  assign \new_Sorter100|14809_  = \new_Sorter100|14708_  | \new_Sorter100|14709_ ;
  assign \new_Sorter100|14810_  = \new_Sorter100|14710_  & \new_Sorter100|14711_ ;
  assign \new_Sorter100|14811_  = \new_Sorter100|14710_  | \new_Sorter100|14711_ ;
  assign \new_Sorter100|14812_  = \new_Sorter100|14712_  & \new_Sorter100|14713_ ;
  assign \new_Sorter100|14813_  = \new_Sorter100|14712_  | \new_Sorter100|14713_ ;
  assign \new_Sorter100|14814_  = \new_Sorter100|14714_  & \new_Sorter100|14715_ ;
  assign \new_Sorter100|14815_  = \new_Sorter100|14714_  | \new_Sorter100|14715_ ;
  assign \new_Sorter100|14816_  = \new_Sorter100|14716_  & \new_Sorter100|14717_ ;
  assign \new_Sorter100|14817_  = \new_Sorter100|14716_  | \new_Sorter100|14717_ ;
  assign \new_Sorter100|14818_  = \new_Sorter100|14718_  & \new_Sorter100|14719_ ;
  assign \new_Sorter100|14819_  = \new_Sorter100|14718_  | \new_Sorter100|14719_ ;
  assign \new_Sorter100|14820_  = \new_Sorter100|14720_  & \new_Sorter100|14721_ ;
  assign \new_Sorter100|14821_  = \new_Sorter100|14720_  | \new_Sorter100|14721_ ;
  assign \new_Sorter100|14822_  = \new_Sorter100|14722_  & \new_Sorter100|14723_ ;
  assign \new_Sorter100|14823_  = \new_Sorter100|14722_  | \new_Sorter100|14723_ ;
  assign \new_Sorter100|14824_  = \new_Sorter100|14724_  & \new_Sorter100|14725_ ;
  assign \new_Sorter100|14825_  = \new_Sorter100|14724_  | \new_Sorter100|14725_ ;
  assign \new_Sorter100|14826_  = \new_Sorter100|14726_  & \new_Sorter100|14727_ ;
  assign \new_Sorter100|14827_  = \new_Sorter100|14726_  | \new_Sorter100|14727_ ;
  assign \new_Sorter100|14828_  = \new_Sorter100|14728_  & \new_Sorter100|14729_ ;
  assign \new_Sorter100|14829_  = \new_Sorter100|14728_  | \new_Sorter100|14729_ ;
  assign \new_Sorter100|14830_  = \new_Sorter100|14730_  & \new_Sorter100|14731_ ;
  assign \new_Sorter100|14831_  = \new_Sorter100|14730_  | \new_Sorter100|14731_ ;
  assign \new_Sorter100|14832_  = \new_Sorter100|14732_  & \new_Sorter100|14733_ ;
  assign \new_Sorter100|14833_  = \new_Sorter100|14732_  | \new_Sorter100|14733_ ;
  assign \new_Sorter100|14834_  = \new_Sorter100|14734_  & \new_Sorter100|14735_ ;
  assign \new_Sorter100|14835_  = \new_Sorter100|14734_  | \new_Sorter100|14735_ ;
  assign \new_Sorter100|14836_  = \new_Sorter100|14736_  & \new_Sorter100|14737_ ;
  assign \new_Sorter100|14837_  = \new_Sorter100|14736_  | \new_Sorter100|14737_ ;
  assign \new_Sorter100|14838_  = \new_Sorter100|14738_  & \new_Sorter100|14739_ ;
  assign \new_Sorter100|14839_  = \new_Sorter100|14738_  | \new_Sorter100|14739_ ;
  assign \new_Sorter100|14840_  = \new_Sorter100|14740_  & \new_Sorter100|14741_ ;
  assign \new_Sorter100|14841_  = \new_Sorter100|14740_  | \new_Sorter100|14741_ ;
  assign \new_Sorter100|14842_  = \new_Sorter100|14742_  & \new_Sorter100|14743_ ;
  assign \new_Sorter100|14843_  = \new_Sorter100|14742_  | \new_Sorter100|14743_ ;
  assign \new_Sorter100|14844_  = \new_Sorter100|14744_  & \new_Sorter100|14745_ ;
  assign \new_Sorter100|14845_  = \new_Sorter100|14744_  | \new_Sorter100|14745_ ;
  assign \new_Sorter100|14846_  = \new_Sorter100|14746_  & \new_Sorter100|14747_ ;
  assign \new_Sorter100|14847_  = \new_Sorter100|14746_  | \new_Sorter100|14747_ ;
  assign \new_Sorter100|14848_  = \new_Sorter100|14748_  & \new_Sorter100|14749_ ;
  assign \new_Sorter100|14849_  = \new_Sorter100|14748_  | \new_Sorter100|14749_ ;
  assign \new_Sorter100|14850_  = \new_Sorter100|14750_  & \new_Sorter100|14751_ ;
  assign \new_Sorter100|14851_  = \new_Sorter100|14750_  | \new_Sorter100|14751_ ;
  assign \new_Sorter100|14852_  = \new_Sorter100|14752_  & \new_Sorter100|14753_ ;
  assign \new_Sorter100|14853_  = \new_Sorter100|14752_  | \new_Sorter100|14753_ ;
  assign \new_Sorter100|14854_  = \new_Sorter100|14754_  & \new_Sorter100|14755_ ;
  assign \new_Sorter100|14855_  = \new_Sorter100|14754_  | \new_Sorter100|14755_ ;
  assign \new_Sorter100|14856_  = \new_Sorter100|14756_  & \new_Sorter100|14757_ ;
  assign \new_Sorter100|14857_  = \new_Sorter100|14756_  | \new_Sorter100|14757_ ;
  assign \new_Sorter100|14858_  = \new_Sorter100|14758_  & \new_Sorter100|14759_ ;
  assign \new_Sorter100|14859_  = \new_Sorter100|14758_  | \new_Sorter100|14759_ ;
  assign \new_Sorter100|14860_  = \new_Sorter100|14760_  & \new_Sorter100|14761_ ;
  assign \new_Sorter100|14861_  = \new_Sorter100|14760_  | \new_Sorter100|14761_ ;
  assign \new_Sorter100|14862_  = \new_Sorter100|14762_  & \new_Sorter100|14763_ ;
  assign \new_Sorter100|14863_  = \new_Sorter100|14762_  | \new_Sorter100|14763_ ;
  assign \new_Sorter100|14864_  = \new_Sorter100|14764_  & \new_Sorter100|14765_ ;
  assign \new_Sorter100|14865_  = \new_Sorter100|14764_  | \new_Sorter100|14765_ ;
  assign \new_Sorter100|14866_  = \new_Sorter100|14766_  & \new_Sorter100|14767_ ;
  assign \new_Sorter100|14867_  = \new_Sorter100|14766_  | \new_Sorter100|14767_ ;
  assign \new_Sorter100|14868_  = \new_Sorter100|14768_  & \new_Sorter100|14769_ ;
  assign \new_Sorter100|14869_  = \new_Sorter100|14768_  | \new_Sorter100|14769_ ;
  assign \new_Sorter100|14870_  = \new_Sorter100|14770_  & \new_Sorter100|14771_ ;
  assign \new_Sorter100|14871_  = \new_Sorter100|14770_  | \new_Sorter100|14771_ ;
  assign \new_Sorter100|14872_  = \new_Sorter100|14772_  & \new_Sorter100|14773_ ;
  assign \new_Sorter100|14873_  = \new_Sorter100|14772_  | \new_Sorter100|14773_ ;
  assign \new_Sorter100|14874_  = \new_Sorter100|14774_  & \new_Sorter100|14775_ ;
  assign \new_Sorter100|14875_  = \new_Sorter100|14774_  | \new_Sorter100|14775_ ;
  assign \new_Sorter100|14876_  = \new_Sorter100|14776_  & \new_Sorter100|14777_ ;
  assign \new_Sorter100|14877_  = \new_Sorter100|14776_  | \new_Sorter100|14777_ ;
  assign \new_Sorter100|14878_  = \new_Sorter100|14778_  & \new_Sorter100|14779_ ;
  assign \new_Sorter100|14879_  = \new_Sorter100|14778_  | \new_Sorter100|14779_ ;
  assign \new_Sorter100|14880_  = \new_Sorter100|14780_  & \new_Sorter100|14781_ ;
  assign \new_Sorter100|14881_  = \new_Sorter100|14780_  | \new_Sorter100|14781_ ;
  assign \new_Sorter100|14882_  = \new_Sorter100|14782_  & \new_Sorter100|14783_ ;
  assign \new_Sorter100|14883_  = \new_Sorter100|14782_  | \new_Sorter100|14783_ ;
  assign \new_Sorter100|14884_  = \new_Sorter100|14784_  & \new_Sorter100|14785_ ;
  assign \new_Sorter100|14885_  = \new_Sorter100|14784_  | \new_Sorter100|14785_ ;
  assign \new_Sorter100|14886_  = \new_Sorter100|14786_  & \new_Sorter100|14787_ ;
  assign \new_Sorter100|14887_  = \new_Sorter100|14786_  | \new_Sorter100|14787_ ;
  assign \new_Sorter100|14888_  = \new_Sorter100|14788_  & \new_Sorter100|14789_ ;
  assign \new_Sorter100|14889_  = \new_Sorter100|14788_  | \new_Sorter100|14789_ ;
  assign \new_Sorter100|14890_  = \new_Sorter100|14790_  & \new_Sorter100|14791_ ;
  assign \new_Sorter100|14891_  = \new_Sorter100|14790_  | \new_Sorter100|14791_ ;
  assign \new_Sorter100|14892_  = \new_Sorter100|14792_  & \new_Sorter100|14793_ ;
  assign \new_Sorter100|14893_  = \new_Sorter100|14792_  | \new_Sorter100|14793_ ;
  assign \new_Sorter100|14894_  = \new_Sorter100|14794_  & \new_Sorter100|14795_ ;
  assign \new_Sorter100|14895_  = \new_Sorter100|14794_  | \new_Sorter100|14795_ ;
  assign \new_Sorter100|14896_  = \new_Sorter100|14796_  & \new_Sorter100|14797_ ;
  assign \new_Sorter100|14897_  = \new_Sorter100|14796_  | \new_Sorter100|14797_ ;
  assign \new_Sorter100|14898_  = \new_Sorter100|14798_  & \new_Sorter100|14799_ ;
  assign \new_Sorter100|14899_  = \new_Sorter100|14798_  | \new_Sorter100|14799_ ;
  assign \new_Sorter100|14900_  = \new_Sorter100|14800_ ;
  assign \new_Sorter100|14999_  = \new_Sorter100|14899_ ;
  assign \new_Sorter100|14901_  = \new_Sorter100|14801_  & \new_Sorter100|14802_ ;
  assign \new_Sorter100|14902_  = \new_Sorter100|14801_  | \new_Sorter100|14802_ ;
  assign \new_Sorter100|14903_  = \new_Sorter100|14803_  & \new_Sorter100|14804_ ;
  assign \new_Sorter100|14904_  = \new_Sorter100|14803_  | \new_Sorter100|14804_ ;
  assign \new_Sorter100|14905_  = \new_Sorter100|14805_  & \new_Sorter100|14806_ ;
  assign \new_Sorter100|14906_  = \new_Sorter100|14805_  | \new_Sorter100|14806_ ;
  assign \new_Sorter100|14907_  = \new_Sorter100|14807_  & \new_Sorter100|14808_ ;
  assign \new_Sorter100|14908_  = \new_Sorter100|14807_  | \new_Sorter100|14808_ ;
  assign \new_Sorter100|14909_  = \new_Sorter100|14809_  & \new_Sorter100|14810_ ;
  assign \new_Sorter100|14910_  = \new_Sorter100|14809_  | \new_Sorter100|14810_ ;
  assign \new_Sorter100|14911_  = \new_Sorter100|14811_  & \new_Sorter100|14812_ ;
  assign \new_Sorter100|14912_  = \new_Sorter100|14811_  | \new_Sorter100|14812_ ;
  assign \new_Sorter100|14913_  = \new_Sorter100|14813_  & \new_Sorter100|14814_ ;
  assign \new_Sorter100|14914_  = \new_Sorter100|14813_  | \new_Sorter100|14814_ ;
  assign \new_Sorter100|14915_  = \new_Sorter100|14815_  & \new_Sorter100|14816_ ;
  assign \new_Sorter100|14916_  = \new_Sorter100|14815_  | \new_Sorter100|14816_ ;
  assign \new_Sorter100|14917_  = \new_Sorter100|14817_  & \new_Sorter100|14818_ ;
  assign \new_Sorter100|14918_  = \new_Sorter100|14817_  | \new_Sorter100|14818_ ;
  assign \new_Sorter100|14919_  = \new_Sorter100|14819_  & \new_Sorter100|14820_ ;
  assign \new_Sorter100|14920_  = \new_Sorter100|14819_  | \new_Sorter100|14820_ ;
  assign \new_Sorter100|14921_  = \new_Sorter100|14821_  & \new_Sorter100|14822_ ;
  assign \new_Sorter100|14922_  = \new_Sorter100|14821_  | \new_Sorter100|14822_ ;
  assign \new_Sorter100|14923_  = \new_Sorter100|14823_  & \new_Sorter100|14824_ ;
  assign \new_Sorter100|14924_  = \new_Sorter100|14823_  | \new_Sorter100|14824_ ;
  assign \new_Sorter100|14925_  = \new_Sorter100|14825_  & \new_Sorter100|14826_ ;
  assign \new_Sorter100|14926_  = \new_Sorter100|14825_  | \new_Sorter100|14826_ ;
  assign \new_Sorter100|14927_  = \new_Sorter100|14827_  & \new_Sorter100|14828_ ;
  assign \new_Sorter100|14928_  = \new_Sorter100|14827_  | \new_Sorter100|14828_ ;
  assign \new_Sorter100|14929_  = \new_Sorter100|14829_  & \new_Sorter100|14830_ ;
  assign \new_Sorter100|14930_  = \new_Sorter100|14829_  | \new_Sorter100|14830_ ;
  assign \new_Sorter100|14931_  = \new_Sorter100|14831_  & \new_Sorter100|14832_ ;
  assign \new_Sorter100|14932_  = \new_Sorter100|14831_  | \new_Sorter100|14832_ ;
  assign \new_Sorter100|14933_  = \new_Sorter100|14833_  & \new_Sorter100|14834_ ;
  assign \new_Sorter100|14934_  = \new_Sorter100|14833_  | \new_Sorter100|14834_ ;
  assign \new_Sorter100|14935_  = \new_Sorter100|14835_  & \new_Sorter100|14836_ ;
  assign \new_Sorter100|14936_  = \new_Sorter100|14835_  | \new_Sorter100|14836_ ;
  assign \new_Sorter100|14937_  = \new_Sorter100|14837_  & \new_Sorter100|14838_ ;
  assign \new_Sorter100|14938_  = \new_Sorter100|14837_  | \new_Sorter100|14838_ ;
  assign \new_Sorter100|14939_  = \new_Sorter100|14839_  & \new_Sorter100|14840_ ;
  assign \new_Sorter100|14940_  = \new_Sorter100|14839_  | \new_Sorter100|14840_ ;
  assign \new_Sorter100|14941_  = \new_Sorter100|14841_  & \new_Sorter100|14842_ ;
  assign \new_Sorter100|14942_  = \new_Sorter100|14841_  | \new_Sorter100|14842_ ;
  assign \new_Sorter100|14943_  = \new_Sorter100|14843_  & \new_Sorter100|14844_ ;
  assign \new_Sorter100|14944_  = \new_Sorter100|14843_  | \new_Sorter100|14844_ ;
  assign \new_Sorter100|14945_  = \new_Sorter100|14845_  & \new_Sorter100|14846_ ;
  assign \new_Sorter100|14946_  = \new_Sorter100|14845_  | \new_Sorter100|14846_ ;
  assign \new_Sorter100|14947_  = \new_Sorter100|14847_  & \new_Sorter100|14848_ ;
  assign \new_Sorter100|14948_  = \new_Sorter100|14847_  | \new_Sorter100|14848_ ;
  assign \new_Sorter100|14949_  = \new_Sorter100|14849_  & \new_Sorter100|14850_ ;
  assign \new_Sorter100|14950_  = \new_Sorter100|14849_  | \new_Sorter100|14850_ ;
  assign \new_Sorter100|14951_  = \new_Sorter100|14851_  & \new_Sorter100|14852_ ;
  assign \new_Sorter100|14952_  = \new_Sorter100|14851_  | \new_Sorter100|14852_ ;
  assign \new_Sorter100|14953_  = \new_Sorter100|14853_  & \new_Sorter100|14854_ ;
  assign \new_Sorter100|14954_  = \new_Sorter100|14853_  | \new_Sorter100|14854_ ;
  assign \new_Sorter100|14955_  = \new_Sorter100|14855_  & \new_Sorter100|14856_ ;
  assign \new_Sorter100|14956_  = \new_Sorter100|14855_  | \new_Sorter100|14856_ ;
  assign \new_Sorter100|14957_  = \new_Sorter100|14857_  & \new_Sorter100|14858_ ;
  assign \new_Sorter100|14958_  = \new_Sorter100|14857_  | \new_Sorter100|14858_ ;
  assign \new_Sorter100|14959_  = \new_Sorter100|14859_  & \new_Sorter100|14860_ ;
  assign \new_Sorter100|14960_  = \new_Sorter100|14859_  | \new_Sorter100|14860_ ;
  assign \new_Sorter100|14961_  = \new_Sorter100|14861_  & \new_Sorter100|14862_ ;
  assign \new_Sorter100|14962_  = \new_Sorter100|14861_  | \new_Sorter100|14862_ ;
  assign \new_Sorter100|14963_  = \new_Sorter100|14863_  & \new_Sorter100|14864_ ;
  assign \new_Sorter100|14964_  = \new_Sorter100|14863_  | \new_Sorter100|14864_ ;
  assign \new_Sorter100|14965_  = \new_Sorter100|14865_  & \new_Sorter100|14866_ ;
  assign \new_Sorter100|14966_  = \new_Sorter100|14865_  | \new_Sorter100|14866_ ;
  assign \new_Sorter100|14967_  = \new_Sorter100|14867_  & \new_Sorter100|14868_ ;
  assign \new_Sorter100|14968_  = \new_Sorter100|14867_  | \new_Sorter100|14868_ ;
  assign \new_Sorter100|14969_  = \new_Sorter100|14869_  & \new_Sorter100|14870_ ;
  assign \new_Sorter100|14970_  = \new_Sorter100|14869_  | \new_Sorter100|14870_ ;
  assign \new_Sorter100|14971_  = \new_Sorter100|14871_  & \new_Sorter100|14872_ ;
  assign \new_Sorter100|14972_  = \new_Sorter100|14871_  | \new_Sorter100|14872_ ;
  assign \new_Sorter100|14973_  = \new_Sorter100|14873_  & \new_Sorter100|14874_ ;
  assign \new_Sorter100|14974_  = \new_Sorter100|14873_  | \new_Sorter100|14874_ ;
  assign \new_Sorter100|14975_  = \new_Sorter100|14875_  & \new_Sorter100|14876_ ;
  assign \new_Sorter100|14976_  = \new_Sorter100|14875_  | \new_Sorter100|14876_ ;
  assign \new_Sorter100|14977_  = \new_Sorter100|14877_  & \new_Sorter100|14878_ ;
  assign \new_Sorter100|14978_  = \new_Sorter100|14877_  | \new_Sorter100|14878_ ;
  assign \new_Sorter100|14979_  = \new_Sorter100|14879_  & \new_Sorter100|14880_ ;
  assign \new_Sorter100|14980_  = \new_Sorter100|14879_  | \new_Sorter100|14880_ ;
  assign \new_Sorter100|14981_  = \new_Sorter100|14881_  & \new_Sorter100|14882_ ;
  assign \new_Sorter100|14982_  = \new_Sorter100|14881_  | \new_Sorter100|14882_ ;
  assign \new_Sorter100|14983_  = \new_Sorter100|14883_  & \new_Sorter100|14884_ ;
  assign \new_Sorter100|14984_  = \new_Sorter100|14883_  | \new_Sorter100|14884_ ;
  assign \new_Sorter100|14985_  = \new_Sorter100|14885_  & \new_Sorter100|14886_ ;
  assign \new_Sorter100|14986_  = \new_Sorter100|14885_  | \new_Sorter100|14886_ ;
  assign \new_Sorter100|14987_  = \new_Sorter100|14887_  & \new_Sorter100|14888_ ;
  assign \new_Sorter100|14988_  = \new_Sorter100|14887_  | \new_Sorter100|14888_ ;
  assign \new_Sorter100|14989_  = \new_Sorter100|14889_  & \new_Sorter100|14890_ ;
  assign \new_Sorter100|14990_  = \new_Sorter100|14889_  | \new_Sorter100|14890_ ;
  assign \new_Sorter100|14991_  = \new_Sorter100|14891_  & \new_Sorter100|14892_ ;
  assign \new_Sorter100|14992_  = \new_Sorter100|14891_  | \new_Sorter100|14892_ ;
  assign \new_Sorter100|14993_  = \new_Sorter100|14893_  & \new_Sorter100|14894_ ;
  assign \new_Sorter100|14994_  = \new_Sorter100|14893_  | \new_Sorter100|14894_ ;
  assign \new_Sorter100|14995_  = \new_Sorter100|14895_  & \new_Sorter100|14896_ ;
  assign \new_Sorter100|14996_  = \new_Sorter100|14895_  | \new_Sorter100|14896_ ;
  assign \new_Sorter100|14997_  = \new_Sorter100|14897_  & \new_Sorter100|14898_ ;
  assign \new_Sorter100|14998_  = \new_Sorter100|14897_  | \new_Sorter100|14898_ ;
  assign \new_Sorter100|15000_  = \new_Sorter100|14900_  & \new_Sorter100|14901_ ;
  assign \new_Sorter100|15001_  = \new_Sorter100|14900_  | \new_Sorter100|14901_ ;
  assign \new_Sorter100|15002_  = \new_Sorter100|14902_  & \new_Sorter100|14903_ ;
  assign \new_Sorter100|15003_  = \new_Sorter100|14902_  | \new_Sorter100|14903_ ;
  assign \new_Sorter100|15004_  = \new_Sorter100|14904_  & \new_Sorter100|14905_ ;
  assign \new_Sorter100|15005_  = \new_Sorter100|14904_  | \new_Sorter100|14905_ ;
  assign \new_Sorter100|15006_  = \new_Sorter100|14906_  & \new_Sorter100|14907_ ;
  assign \new_Sorter100|15007_  = \new_Sorter100|14906_  | \new_Sorter100|14907_ ;
  assign \new_Sorter100|15008_  = \new_Sorter100|14908_  & \new_Sorter100|14909_ ;
  assign \new_Sorter100|15009_  = \new_Sorter100|14908_  | \new_Sorter100|14909_ ;
  assign \new_Sorter100|15010_  = \new_Sorter100|14910_  & \new_Sorter100|14911_ ;
  assign \new_Sorter100|15011_  = \new_Sorter100|14910_  | \new_Sorter100|14911_ ;
  assign \new_Sorter100|15012_  = \new_Sorter100|14912_  & \new_Sorter100|14913_ ;
  assign \new_Sorter100|15013_  = \new_Sorter100|14912_  | \new_Sorter100|14913_ ;
  assign \new_Sorter100|15014_  = \new_Sorter100|14914_  & \new_Sorter100|14915_ ;
  assign \new_Sorter100|15015_  = \new_Sorter100|14914_  | \new_Sorter100|14915_ ;
  assign \new_Sorter100|15016_  = \new_Sorter100|14916_  & \new_Sorter100|14917_ ;
  assign \new_Sorter100|15017_  = \new_Sorter100|14916_  | \new_Sorter100|14917_ ;
  assign \new_Sorter100|15018_  = \new_Sorter100|14918_  & \new_Sorter100|14919_ ;
  assign \new_Sorter100|15019_  = \new_Sorter100|14918_  | \new_Sorter100|14919_ ;
  assign \new_Sorter100|15020_  = \new_Sorter100|14920_  & \new_Sorter100|14921_ ;
  assign \new_Sorter100|15021_  = \new_Sorter100|14920_  | \new_Sorter100|14921_ ;
  assign \new_Sorter100|15022_  = \new_Sorter100|14922_  & \new_Sorter100|14923_ ;
  assign \new_Sorter100|15023_  = \new_Sorter100|14922_  | \new_Sorter100|14923_ ;
  assign \new_Sorter100|15024_  = \new_Sorter100|14924_  & \new_Sorter100|14925_ ;
  assign \new_Sorter100|15025_  = \new_Sorter100|14924_  | \new_Sorter100|14925_ ;
  assign \new_Sorter100|15026_  = \new_Sorter100|14926_  & \new_Sorter100|14927_ ;
  assign \new_Sorter100|15027_  = \new_Sorter100|14926_  | \new_Sorter100|14927_ ;
  assign \new_Sorter100|15028_  = \new_Sorter100|14928_  & \new_Sorter100|14929_ ;
  assign \new_Sorter100|15029_  = \new_Sorter100|14928_  | \new_Sorter100|14929_ ;
  assign \new_Sorter100|15030_  = \new_Sorter100|14930_  & \new_Sorter100|14931_ ;
  assign \new_Sorter100|15031_  = \new_Sorter100|14930_  | \new_Sorter100|14931_ ;
  assign \new_Sorter100|15032_  = \new_Sorter100|14932_  & \new_Sorter100|14933_ ;
  assign \new_Sorter100|15033_  = \new_Sorter100|14932_  | \new_Sorter100|14933_ ;
  assign \new_Sorter100|15034_  = \new_Sorter100|14934_  & \new_Sorter100|14935_ ;
  assign \new_Sorter100|15035_  = \new_Sorter100|14934_  | \new_Sorter100|14935_ ;
  assign \new_Sorter100|15036_  = \new_Sorter100|14936_  & \new_Sorter100|14937_ ;
  assign \new_Sorter100|15037_  = \new_Sorter100|14936_  | \new_Sorter100|14937_ ;
  assign \new_Sorter100|15038_  = \new_Sorter100|14938_  & \new_Sorter100|14939_ ;
  assign \new_Sorter100|15039_  = \new_Sorter100|14938_  | \new_Sorter100|14939_ ;
  assign \new_Sorter100|15040_  = \new_Sorter100|14940_  & \new_Sorter100|14941_ ;
  assign \new_Sorter100|15041_  = \new_Sorter100|14940_  | \new_Sorter100|14941_ ;
  assign \new_Sorter100|15042_  = \new_Sorter100|14942_  & \new_Sorter100|14943_ ;
  assign \new_Sorter100|15043_  = \new_Sorter100|14942_  | \new_Sorter100|14943_ ;
  assign \new_Sorter100|15044_  = \new_Sorter100|14944_  & \new_Sorter100|14945_ ;
  assign \new_Sorter100|15045_  = \new_Sorter100|14944_  | \new_Sorter100|14945_ ;
  assign \new_Sorter100|15046_  = \new_Sorter100|14946_  & \new_Sorter100|14947_ ;
  assign \new_Sorter100|15047_  = \new_Sorter100|14946_  | \new_Sorter100|14947_ ;
  assign \new_Sorter100|15048_  = \new_Sorter100|14948_  & \new_Sorter100|14949_ ;
  assign \new_Sorter100|15049_  = \new_Sorter100|14948_  | \new_Sorter100|14949_ ;
  assign \new_Sorter100|15050_  = \new_Sorter100|14950_  & \new_Sorter100|14951_ ;
  assign \new_Sorter100|15051_  = \new_Sorter100|14950_  | \new_Sorter100|14951_ ;
  assign \new_Sorter100|15052_  = \new_Sorter100|14952_  & \new_Sorter100|14953_ ;
  assign \new_Sorter100|15053_  = \new_Sorter100|14952_  | \new_Sorter100|14953_ ;
  assign \new_Sorter100|15054_  = \new_Sorter100|14954_  & \new_Sorter100|14955_ ;
  assign \new_Sorter100|15055_  = \new_Sorter100|14954_  | \new_Sorter100|14955_ ;
  assign \new_Sorter100|15056_  = \new_Sorter100|14956_  & \new_Sorter100|14957_ ;
  assign \new_Sorter100|15057_  = \new_Sorter100|14956_  | \new_Sorter100|14957_ ;
  assign \new_Sorter100|15058_  = \new_Sorter100|14958_  & \new_Sorter100|14959_ ;
  assign \new_Sorter100|15059_  = \new_Sorter100|14958_  | \new_Sorter100|14959_ ;
  assign \new_Sorter100|15060_  = \new_Sorter100|14960_  & \new_Sorter100|14961_ ;
  assign \new_Sorter100|15061_  = \new_Sorter100|14960_  | \new_Sorter100|14961_ ;
  assign \new_Sorter100|15062_  = \new_Sorter100|14962_  & \new_Sorter100|14963_ ;
  assign \new_Sorter100|15063_  = \new_Sorter100|14962_  | \new_Sorter100|14963_ ;
  assign \new_Sorter100|15064_  = \new_Sorter100|14964_  & \new_Sorter100|14965_ ;
  assign \new_Sorter100|15065_  = \new_Sorter100|14964_  | \new_Sorter100|14965_ ;
  assign \new_Sorter100|15066_  = \new_Sorter100|14966_  & \new_Sorter100|14967_ ;
  assign \new_Sorter100|15067_  = \new_Sorter100|14966_  | \new_Sorter100|14967_ ;
  assign \new_Sorter100|15068_  = \new_Sorter100|14968_  & \new_Sorter100|14969_ ;
  assign \new_Sorter100|15069_  = \new_Sorter100|14968_  | \new_Sorter100|14969_ ;
  assign \new_Sorter100|15070_  = \new_Sorter100|14970_  & \new_Sorter100|14971_ ;
  assign \new_Sorter100|15071_  = \new_Sorter100|14970_  | \new_Sorter100|14971_ ;
  assign \new_Sorter100|15072_  = \new_Sorter100|14972_  & \new_Sorter100|14973_ ;
  assign \new_Sorter100|15073_  = \new_Sorter100|14972_  | \new_Sorter100|14973_ ;
  assign \new_Sorter100|15074_  = \new_Sorter100|14974_  & \new_Sorter100|14975_ ;
  assign \new_Sorter100|15075_  = \new_Sorter100|14974_  | \new_Sorter100|14975_ ;
  assign \new_Sorter100|15076_  = \new_Sorter100|14976_  & \new_Sorter100|14977_ ;
  assign \new_Sorter100|15077_  = \new_Sorter100|14976_  | \new_Sorter100|14977_ ;
  assign \new_Sorter100|15078_  = \new_Sorter100|14978_  & \new_Sorter100|14979_ ;
  assign \new_Sorter100|15079_  = \new_Sorter100|14978_  | \new_Sorter100|14979_ ;
  assign \new_Sorter100|15080_  = \new_Sorter100|14980_  & \new_Sorter100|14981_ ;
  assign \new_Sorter100|15081_  = \new_Sorter100|14980_  | \new_Sorter100|14981_ ;
  assign \new_Sorter100|15082_  = \new_Sorter100|14982_  & \new_Sorter100|14983_ ;
  assign \new_Sorter100|15083_  = \new_Sorter100|14982_  | \new_Sorter100|14983_ ;
  assign \new_Sorter100|15084_  = \new_Sorter100|14984_  & \new_Sorter100|14985_ ;
  assign \new_Sorter100|15085_  = \new_Sorter100|14984_  | \new_Sorter100|14985_ ;
  assign \new_Sorter100|15086_  = \new_Sorter100|14986_  & \new_Sorter100|14987_ ;
  assign \new_Sorter100|15087_  = \new_Sorter100|14986_  | \new_Sorter100|14987_ ;
  assign \new_Sorter100|15088_  = \new_Sorter100|14988_  & \new_Sorter100|14989_ ;
  assign \new_Sorter100|15089_  = \new_Sorter100|14988_  | \new_Sorter100|14989_ ;
  assign \new_Sorter100|15090_  = \new_Sorter100|14990_  & \new_Sorter100|14991_ ;
  assign \new_Sorter100|15091_  = \new_Sorter100|14990_  | \new_Sorter100|14991_ ;
  assign \new_Sorter100|15092_  = \new_Sorter100|14992_  & \new_Sorter100|14993_ ;
  assign \new_Sorter100|15093_  = \new_Sorter100|14992_  | \new_Sorter100|14993_ ;
  assign \new_Sorter100|15094_  = \new_Sorter100|14994_  & \new_Sorter100|14995_ ;
  assign \new_Sorter100|15095_  = \new_Sorter100|14994_  | \new_Sorter100|14995_ ;
  assign \new_Sorter100|15096_  = \new_Sorter100|14996_  & \new_Sorter100|14997_ ;
  assign \new_Sorter100|15097_  = \new_Sorter100|14996_  | \new_Sorter100|14997_ ;
  assign \new_Sorter100|15098_  = \new_Sorter100|14998_  & \new_Sorter100|14999_ ;
  assign \new_Sorter100|15099_  = \new_Sorter100|14998_  | \new_Sorter100|14999_ ;
  assign \new_Sorter100|15100_  = \new_Sorter100|15000_ ;
  assign \new_Sorter100|15199_  = \new_Sorter100|15099_ ;
  assign \new_Sorter100|15101_  = \new_Sorter100|15001_  & \new_Sorter100|15002_ ;
  assign \new_Sorter100|15102_  = \new_Sorter100|15001_  | \new_Sorter100|15002_ ;
  assign \new_Sorter100|15103_  = \new_Sorter100|15003_  & \new_Sorter100|15004_ ;
  assign \new_Sorter100|15104_  = \new_Sorter100|15003_  | \new_Sorter100|15004_ ;
  assign \new_Sorter100|15105_  = \new_Sorter100|15005_  & \new_Sorter100|15006_ ;
  assign \new_Sorter100|15106_  = \new_Sorter100|15005_  | \new_Sorter100|15006_ ;
  assign \new_Sorter100|15107_  = \new_Sorter100|15007_  & \new_Sorter100|15008_ ;
  assign \new_Sorter100|15108_  = \new_Sorter100|15007_  | \new_Sorter100|15008_ ;
  assign \new_Sorter100|15109_  = \new_Sorter100|15009_  & \new_Sorter100|15010_ ;
  assign \new_Sorter100|15110_  = \new_Sorter100|15009_  | \new_Sorter100|15010_ ;
  assign \new_Sorter100|15111_  = \new_Sorter100|15011_  & \new_Sorter100|15012_ ;
  assign \new_Sorter100|15112_  = \new_Sorter100|15011_  | \new_Sorter100|15012_ ;
  assign \new_Sorter100|15113_  = \new_Sorter100|15013_  & \new_Sorter100|15014_ ;
  assign \new_Sorter100|15114_  = \new_Sorter100|15013_  | \new_Sorter100|15014_ ;
  assign \new_Sorter100|15115_  = \new_Sorter100|15015_  & \new_Sorter100|15016_ ;
  assign \new_Sorter100|15116_  = \new_Sorter100|15015_  | \new_Sorter100|15016_ ;
  assign \new_Sorter100|15117_  = \new_Sorter100|15017_  & \new_Sorter100|15018_ ;
  assign \new_Sorter100|15118_  = \new_Sorter100|15017_  | \new_Sorter100|15018_ ;
  assign \new_Sorter100|15119_  = \new_Sorter100|15019_  & \new_Sorter100|15020_ ;
  assign \new_Sorter100|15120_  = \new_Sorter100|15019_  | \new_Sorter100|15020_ ;
  assign \new_Sorter100|15121_  = \new_Sorter100|15021_  & \new_Sorter100|15022_ ;
  assign \new_Sorter100|15122_  = \new_Sorter100|15021_  | \new_Sorter100|15022_ ;
  assign \new_Sorter100|15123_  = \new_Sorter100|15023_  & \new_Sorter100|15024_ ;
  assign \new_Sorter100|15124_  = \new_Sorter100|15023_  | \new_Sorter100|15024_ ;
  assign \new_Sorter100|15125_  = \new_Sorter100|15025_  & \new_Sorter100|15026_ ;
  assign \new_Sorter100|15126_  = \new_Sorter100|15025_  | \new_Sorter100|15026_ ;
  assign \new_Sorter100|15127_  = \new_Sorter100|15027_  & \new_Sorter100|15028_ ;
  assign \new_Sorter100|15128_  = \new_Sorter100|15027_  | \new_Sorter100|15028_ ;
  assign \new_Sorter100|15129_  = \new_Sorter100|15029_  & \new_Sorter100|15030_ ;
  assign \new_Sorter100|15130_  = \new_Sorter100|15029_  | \new_Sorter100|15030_ ;
  assign \new_Sorter100|15131_  = \new_Sorter100|15031_  & \new_Sorter100|15032_ ;
  assign \new_Sorter100|15132_  = \new_Sorter100|15031_  | \new_Sorter100|15032_ ;
  assign \new_Sorter100|15133_  = \new_Sorter100|15033_  & \new_Sorter100|15034_ ;
  assign \new_Sorter100|15134_  = \new_Sorter100|15033_  | \new_Sorter100|15034_ ;
  assign \new_Sorter100|15135_  = \new_Sorter100|15035_  & \new_Sorter100|15036_ ;
  assign \new_Sorter100|15136_  = \new_Sorter100|15035_  | \new_Sorter100|15036_ ;
  assign \new_Sorter100|15137_  = \new_Sorter100|15037_  & \new_Sorter100|15038_ ;
  assign \new_Sorter100|15138_  = \new_Sorter100|15037_  | \new_Sorter100|15038_ ;
  assign \new_Sorter100|15139_  = \new_Sorter100|15039_  & \new_Sorter100|15040_ ;
  assign \new_Sorter100|15140_  = \new_Sorter100|15039_  | \new_Sorter100|15040_ ;
  assign \new_Sorter100|15141_  = \new_Sorter100|15041_  & \new_Sorter100|15042_ ;
  assign \new_Sorter100|15142_  = \new_Sorter100|15041_  | \new_Sorter100|15042_ ;
  assign \new_Sorter100|15143_  = \new_Sorter100|15043_  & \new_Sorter100|15044_ ;
  assign \new_Sorter100|15144_  = \new_Sorter100|15043_  | \new_Sorter100|15044_ ;
  assign \new_Sorter100|15145_  = \new_Sorter100|15045_  & \new_Sorter100|15046_ ;
  assign \new_Sorter100|15146_  = \new_Sorter100|15045_  | \new_Sorter100|15046_ ;
  assign \new_Sorter100|15147_  = \new_Sorter100|15047_  & \new_Sorter100|15048_ ;
  assign \new_Sorter100|15148_  = \new_Sorter100|15047_  | \new_Sorter100|15048_ ;
  assign \new_Sorter100|15149_  = \new_Sorter100|15049_  & \new_Sorter100|15050_ ;
  assign \new_Sorter100|15150_  = \new_Sorter100|15049_  | \new_Sorter100|15050_ ;
  assign \new_Sorter100|15151_  = \new_Sorter100|15051_  & \new_Sorter100|15052_ ;
  assign \new_Sorter100|15152_  = \new_Sorter100|15051_  | \new_Sorter100|15052_ ;
  assign \new_Sorter100|15153_  = \new_Sorter100|15053_  & \new_Sorter100|15054_ ;
  assign \new_Sorter100|15154_  = \new_Sorter100|15053_  | \new_Sorter100|15054_ ;
  assign \new_Sorter100|15155_  = \new_Sorter100|15055_  & \new_Sorter100|15056_ ;
  assign \new_Sorter100|15156_  = \new_Sorter100|15055_  | \new_Sorter100|15056_ ;
  assign \new_Sorter100|15157_  = \new_Sorter100|15057_  & \new_Sorter100|15058_ ;
  assign \new_Sorter100|15158_  = \new_Sorter100|15057_  | \new_Sorter100|15058_ ;
  assign \new_Sorter100|15159_  = \new_Sorter100|15059_  & \new_Sorter100|15060_ ;
  assign \new_Sorter100|15160_  = \new_Sorter100|15059_  | \new_Sorter100|15060_ ;
  assign \new_Sorter100|15161_  = \new_Sorter100|15061_  & \new_Sorter100|15062_ ;
  assign \new_Sorter100|15162_  = \new_Sorter100|15061_  | \new_Sorter100|15062_ ;
  assign \new_Sorter100|15163_  = \new_Sorter100|15063_  & \new_Sorter100|15064_ ;
  assign \new_Sorter100|15164_  = \new_Sorter100|15063_  | \new_Sorter100|15064_ ;
  assign \new_Sorter100|15165_  = \new_Sorter100|15065_  & \new_Sorter100|15066_ ;
  assign \new_Sorter100|15166_  = \new_Sorter100|15065_  | \new_Sorter100|15066_ ;
  assign \new_Sorter100|15167_  = \new_Sorter100|15067_  & \new_Sorter100|15068_ ;
  assign \new_Sorter100|15168_  = \new_Sorter100|15067_  | \new_Sorter100|15068_ ;
  assign \new_Sorter100|15169_  = \new_Sorter100|15069_  & \new_Sorter100|15070_ ;
  assign \new_Sorter100|15170_  = \new_Sorter100|15069_  | \new_Sorter100|15070_ ;
  assign \new_Sorter100|15171_  = \new_Sorter100|15071_  & \new_Sorter100|15072_ ;
  assign \new_Sorter100|15172_  = \new_Sorter100|15071_  | \new_Sorter100|15072_ ;
  assign \new_Sorter100|15173_  = \new_Sorter100|15073_  & \new_Sorter100|15074_ ;
  assign \new_Sorter100|15174_  = \new_Sorter100|15073_  | \new_Sorter100|15074_ ;
  assign \new_Sorter100|15175_  = \new_Sorter100|15075_  & \new_Sorter100|15076_ ;
  assign \new_Sorter100|15176_  = \new_Sorter100|15075_  | \new_Sorter100|15076_ ;
  assign \new_Sorter100|15177_  = \new_Sorter100|15077_  & \new_Sorter100|15078_ ;
  assign \new_Sorter100|15178_  = \new_Sorter100|15077_  | \new_Sorter100|15078_ ;
  assign \new_Sorter100|15179_  = \new_Sorter100|15079_  & \new_Sorter100|15080_ ;
  assign \new_Sorter100|15180_  = \new_Sorter100|15079_  | \new_Sorter100|15080_ ;
  assign \new_Sorter100|15181_  = \new_Sorter100|15081_  & \new_Sorter100|15082_ ;
  assign \new_Sorter100|15182_  = \new_Sorter100|15081_  | \new_Sorter100|15082_ ;
  assign \new_Sorter100|15183_  = \new_Sorter100|15083_  & \new_Sorter100|15084_ ;
  assign \new_Sorter100|15184_  = \new_Sorter100|15083_  | \new_Sorter100|15084_ ;
  assign \new_Sorter100|15185_  = \new_Sorter100|15085_  & \new_Sorter100|15086_ ;
  assign \new_Sorter100|15186_  = \new_Sorter100|15085_  | \new_Sorter100|15086_ ;
  assign \new_Sorter100|15187_  = \new_Sorter100|15087_  & \new_Sorter100|15088_ ;
  assign \new_Sorter100|15188_  = \new_Sorter100|15087_  | \new_Sorter100|15088_ ;
  assign \new_Sorter100|15189_  = \new_Sorter100|15089_  & \new_Sorter100|15090_ ;
  assign \new_Sorter100|15190_  = \new_Sorter100|15089_  | \new_Sorter100|15090_ ;
  assign \new_Sorter100|15191_  = \new_Sorter100|15091_  & \new_Sorter100|15092_ ;
  assign \new_Sorter100|15192_  = \new_Sorter100|15091_  | \new_Sorter100|15092_ ;
  assign \new_Sorter100|15193_  = \new_Sorter100|15093_  & \new_Sorter100|15094_ ;
  assign \new_Sorter100|15194_  = \new_Sorter100|15093_  | \new_Sorter100|15094_ ;
  assign \new_Sorter100|15195_  = \new_Sorter100|15095_  & \new_Sorter100|15096_ ;
  assign \new_Sorter100|15196_  = \new_Sorter100|15095_  | \new_Sorter100|15096_ ;
  assign \new_Sorter100|15197_  = \new_Sorter100|15097_  & \new_Sorter100|15098_ ;
  assign \new_Sorter100|15198_  = \new_Sorter100|15097_  | \new_Sorter100|15098_ ;
  assign \new_Sorter100|15200_  = \new_Sorter100|15100_  & \new_Sorter100|15101_ ;
  assign \new_Sorter100|15201_  = \new_Sorter100|15100_  | \new_Sorter100|15101_ ;
  assign \new_Sorter100|15202_  = \new_Sorter100|15102_  & \new_Sorter100|15103_ ;
  assign \new_Sorter100|15203_  = \new_Sorter100|15102_  | \new_Sorter100|15103_ ;
  assign \new_Sorter100|15204_  = \new_Sorter100|15104_  & \new_Sorter100|15105_ ;
  assign \new_Sorter100|15205_  = \new_Sorter100|15104_  | \new_Sorter100|15105_ ;
  assign \new_Sorter100|15206_  = \new_Sorter100|15106_  & \new_Sorter100|15107_ ;
  assign \new_Sorter100|15207_  = \new_Sorter100|15106_  | \new_Sorter100|15107_ ;
  assign \new_Sorter100|15208_  = \new_Sorter100|15108_  & \new_Sorter100|15109_ ;
  assign \new_Sorter100|15209_  = \new_Sorter100|15108_  | \new_Sorter100|15109_ ;
  assign \new_Sorter100|15210_  = \new_Sorter100|15110_  & \new_Sorter100|15111_ ;
  assign \new_Sorter100|15211_  = \new_Sorter100|15110_  | \new_Sorter100|15111_ ;
  assign \new_Sorter100|15212_  = \new_Sorter100|15112_  & \new_Sorter100|15113_ ;
  assign \new_Sorter100|15213_  = \new_Sorter100|15112_  | \new_Sorter100|15113_ ;
  assign \new_Sorter100|15214_  = \new_Sorter100|15114_  & \new_Sorter100|15115_ ;
  assign \new_Sorter100|15215_  = \new_Sorter100|15114_  | \new_Sorter100|15115_ ;
  assign \new_Sorter100|15216_  = \new_Sorter100|15116_  & \new_Sorter100|15117_ ;
  assign \new_Sorter100|15217_  = \new_Sorter100|15116_  | \new_Sorter100|15117_ ;
  assign \new_Sorter100|15218_  = \new_Sorter100|15118_  & \new_Sorter100|15119_ ;
  assign \new_Sorter100|15219_  = \new_Sorter100|15118_  | \new_Sorter100|15119_ ;
  assign \new_Sorter100|15220_  = \new_Sorter100|15120_  & \new_Sorter100|15121_ ;
  assign \new_Sorter100|15221_  = \new_Sorter100|15120_  | \new_Sorter100|15121_ ;
  assign \new_Sorter100|15222_  = \new_Sorter100|15122_  & \new_Sorter100|15123_ ;
  assign \new_Sorter100|15223_  = \new_Sorter100|15122_  | \new_Sorter100|15123_ ;
  assign \new_Sorter100|15224_  = \new_Sorter100|15124_  & \new_Sorter100|15125_ ;
  assign \new_Sorter100|15225_  = \new_Sorter100|15124_  | \new_Sorter100|15125_ ;
  assign \new_Sorter100|15226_  = \new_Sorter100|15126_  & \new_Sorter100|15127_ ;
  assign \new_Sorter100|15227_  = \new_Sorter100|15126_  | \new_Sorter100|15127_ ;
  assign \new_Sorter100|15228_  = \new_Sorter100|15128_  & \new_Sorter100|15129_ ;
  assign \new_Sorter100|15229_  = \new_Sorter100|15128_  | \new_Sorter100|15129_ ;
  assign \new_Sorter100|15230_  = \new_Sorter100|15130_  & \new_Sorter100|15131_ ;
  assign \new_Sorter100|15231_  = \new_Sorter100|15130_  | \new_Sorter100|15131_ ;
  assign \new_Sorter100|15232_  = \new_Sorter100|15132_  & \new_Sorter100|15133_ ;
  assign \new_Sorter100|15233_  = \new_Sorter100|15132_  | \new_Sorter100|15133_ ;
  assign \new_Sorter100|15234_  = \new_Sorter100|15134_  & \new_Sorter100|15135_ ;
  assign \new_Sorter100|15235_  = \new_Sorter100|15134_  | \new_Sorter100|15135_ ;
  assign \new_Sorter100|15236_  = \new_Sorter100|15136_  & \new_Sorter100|15137_ ;
  assign \new_Sorter100|15237_  = \new_Sorter100|15136_  | \new_Sorter100|15137_ ;
  assign \new_Sorter100|15238_  = \new_Sorter100|15138_  & \new_Sorter100|15139_ ;
  assign \new_Sorter100|15239_  = \new_Sorter100|15138_  | \new_Sorter100|15139_ ;
  assign \new_Sorter100|15240_  = \new_Sorter100|15140_  & \new_Sorter100|15141_ ;
  assign \new_Sorter100|15241_  = \new_Sorter100|15140_  | \new_Sorter100|15141_ ;
  assign \new_Sorter100|15242_  = \new_Sorter100|15142_  & \new_Sorter100|15143_ ;
  assign \new_Sorter100|15243_  = \new_Sorter100|15142_  | \new_Sorter100|15143_ ;
  assign \new_Sorter100|15244_  = \new_Sorter100|15144_  & \new_Sorter100|15145_ ;
  assign \new_Sorter100|15245_  = \new_Sorter100|15144_  | \new_Sorter100|15145_ ;
  assign \new_Sorter100|15246_  = \new_Sorter100|15146_  & \new_Sorter100|15147_ ;
  assign \new_Sorter100|15247_  = \new_Sorter100|15146_  | \new_Sorter100|15147_ ;
  assign \new_Sorter100|15248_  = \new_Sorter100|15148_  & \new_Sorter100|15149_ ;
  assign \new_Sorter100|15249_  = \new_Sorter100|15148_  | \new_Sorter100|15149_ ;
  assign \new_Sorter100|15250_  = \new_Sorter100|15150_  & \new_Sorter100|15151_ ;
  assign \new_Sorter100|15251_  = \new_Sorter100|15150_  | \new_Sorter100|15151_ ;
  assign \new_Sorter100|15252_  = \new_Sorter100|15152_  & \new_Sorter100|15153_ ;
  assign \new_Sorter100|15253_  = \new_Sorter100|15152_  | \new_Sorter100|15153_ ;
  assign \new_Sorter100|15254_  = \new_Sorter100|15154_  & \new_Sorter100|15155_ ;
  assign \new_Sorter100|15255_  = \new_Sorter100|15154_  | \new_Sorter100|15155_ ;
  assign \new_Sorter100|15256_  = \new_Sorter100|15156_  & \new_Sorter100|15157_ ;
  assign \new_Sorter100|15257_  = \new_Sorter100|15156_  | \new_Sorter100|15157_ ;
  assign \new_Sorter100|15258_  = \new_Sorter100|15158_  & \new_Sorter100|15159_ ;
  assign \new_Sorter100|15259_  = \new_Sorter100|15158_  | \new_Sorter100|15159_ ;
  assign \new_Sorter100|15260_  = \new_Sorter100|15160_  & \new_Sorter100|15161_ ;
  assign \new_Sorter100|15261_  = \new_Sorter100|15160_  | \new_Sorter100|15161_ ;
  assign \new_Sorter100|15262_  = \new_Sorter100|15162_  & \new_Sorter100|15163_ ;
  assign \new_Sorter100|15263_  = \new_Sorter100|15162_  | \new_Sorter100|15163_ ;
  assign \new_Sorter100|15264_  = \new_Sorter100|15164_  & \new_Sorter100|15165_ ;
  assign \new_Sorter100|15265_  = \new_Sorter100|15164_  | \new_Sorter100|15165_ ;
  assign \new_Sorter100|15266_  = \new_Sorter100|15166_  & \new_Sorter100|15167_ ;
  assign \new_Sorter100|15267_  = \new_Sorter100|15166_  | \new_Sorter100|15167_ ;
  assign \new_Sorter100|15268_  = \new_Sorter100|15168_  & \new_Sorter100|15169_ ;
  assign \new_Sorter100|15269_  = \new_Sorter100|15168_  | \new_Sorter100|15169_ ;
  assign \new_Sorter100|15270_  = \new_Sorter100|15170_  & \new_Sorter100|15171_ ;
  assign \new_Sorter100|15271_  = \new_Sorter100|15170_  | \new_Sorter100|15171_ ;
  assign \new_Sorter100|15272_  = \new_Sorter100|15172_  & \new_Sorter100|15173_ ;
  assign \new_Sorter100|15273_  = \new_Sorter100|15172_  | \new_Sorter100|15173_ ;
  assign \new_Sorter100|15274_  = \new_Sorter100|15174_  & \new_Sorter100|15175_ ;
  assign \new_Sorter100|15275_  = \new_Sorter100|15174_  | \new_Sorter100|15175_ ;
  assign \new_Sorter100|15276_  = \new_Sorter100|15176_  & \new_Sorter100|15177_ ;
  assign \new_Sorter100|15277_  = \new_Sorter100|15176_  | \new_Sorter100|15177_ ;
  assign \new_Sorter100|15278_  = \new_Sorter100|15178_  & \new_Sorter100|15179_ ;
  assign \new_Sorter100|15279_  = \new_Sorter100|15178_  | \new_Sorter100|15179_ ;
  assign \new_Sorter100|15280_  = \new_Sorter100|15180_  & \new_Sorter100|15181_ ;
  assign \new_Sorter100|15281_  = \new_Sorter100|15180_  | \new_Sorter100|15181_ ;
  assign \new_Sorter100|15282_  = \new_Sorter100|15182_  & \new_Sorter100|15183_ ;
  assign \new_Sorter100|15283_  = \new_Sorter100|15182_  | \new_Sorter100|15183_ ;
  assign \new_Sorter100|15284_  = \new_Sorter100|15184_  & \new_Sorter100|15185_ ;
  assign \new_Sorter100|15285_  = \new_Sorter100|15184_  | \new_Sorter100|15185_ ;
  assign \new_Sorter100|15286_  = \new_Sorter100|15186_  & \new_Sorter100|15187_ ;
  assign \new_Sorter100|15287_  = \new_Sorter100|15186_  | \new_Sorter100|15187_ ;
  assign \new_Sorter100|15288_  = \new_Sorter100|15188_  & \new_Sorter100|15189_ ;
  assign \new_Sorter100|15289_  = \new_Sorter100|15188_  | \new_Sorter100|15189_ ;
  assign \new_Sorter100|15290_  = \new_Sorter100|15190_  & \new_Sorter100|15191_ ;
  assign \new_Sorter100|15291_  = \new_Sorter100|15190_  | \new_Sorter100|15191_ ;
  assign \new_Sorter100|15292_  = \new_Sorter100|15192_  & \new_Sorter100|15193_ ;
  assign \new_Sorter100|15293_  = \new_Sorter100|15192_  | \new_Sorter100|15193_ ;
  assign \new_Sorter100|15294_  = \new_Sorter100|15194_  & \new_Sorter100|15195_ ;
  assign \new_Sorter100|15295_  = \new_Sorter100|15194_  | \new_Sorter100|15195_ ;
  assign \new_Sorter100|15296_  = \new_Sorter100|15196_  & \new_Sorter100|15197_ ;
  assign \new_Sorter100|15297_  = \new_Sorter100|15196_  | \new_Sorter100|15197_ ;
  assign \new_Sorter100|15298_  = \new_Sorter100|15198_  & \new_Sorter100|15199_ ;
  assign \new_Sorter100|15299_  = \new_Sorter100|15198_  | \new_Sorter100|15199_ ;
  assign \new_Sorter100|15300_  = \new_Sorter100|15200_ ;
  assign \new_Sorter100|15399_  = \new_Sorter100|15299_ ;
  assign \new_Sorter100|15301_  = \new_Sorter100|15201_  & \new_Sorter100|15202_ ;
  assign \new_Sorter100|15302_  = \new_Sorter100|15201_  | \new_Sorter100|15202_ ;
  assign \new_Sorter100|15303_  = \new_Sorter100|15203_  & \new_Sorter100|15204_ ;
  assign \new_Sorter100|15304_  = \new_Sorter100|15203_  | \new_Sorter100|15204_ ;
  assign \new_Sorter100|15305_  = \new_Sorter100|15205_  & \new_Sorter100|15206_ ;
  assign \new_Sorter100|15306_  = \new_Sorter100|15205_  | \new_Sorter100|15206_ ;
  assign \new_Sorter100|15307_  = \new_Sorter100|15207_  & \new_Sorter100|15208_ ;
  assign \new_Sorter100|15308_  = \new_Sorter100|15207_  | \new_Sorter100|15208_ ;
  assign \new_Sorter100|15309_  = \new_Sorter100|15209_  & \new_Sorter100|15210_ ;
  assign \new_Sorter100|15310_  = \new_Sorter100|15209_  | \new_Sorter100|15210_ ;
  assign \new_Sorter100|15311_  = \new_Sorter100|15211_  & \new_Sorter100|15212_ ;
  assign \new_Sorter100|15312_  = \new_Sorter100|15211_  | \new_Sorter100|15212_ ;
  assign \new_Sorter100|15313_  = \new_Sorter100|15213_  & \new_Sorter100|15214_ ;
  assign \new_Sorter100|15314_  = \new_Sorter100|15213_  | \new_Sorter100|15214_ ;
  assign \new_Sorter100|15315_  = \new_Sorter100|15215_  & \new_Sorter100|15216_ ;
  assign \new_Sorter100|15316_  = \new_Sorter100|15215_  | \new_Sorter100|15216_ ;
  assign \new_Sorter100|15317_  = \new_Sorter100|15217_  & \new_Sorter100|15218_ ;
  assign \new_Sorter100|15318_  = \new_Sorter100|15217_  | \new_Sorter100|15218_ ;
  assign \new_Sorter100|15319_  = \new_Sorter100|15219_  & \new_Sorter100|15220_ ;
  assign \new_Sorter100|15320_  = \new_Sorter100|15219_  | \new_Sorter100|15220_ ;
  assign \new_Sorter100|15321_  = \new_Sorter100|15221_  & \new_Sorter100|15222_ ;
  assign \new_Sorter100|15322_  = \new_Sorter100|15221_  | \new_Sorter100|15222_ ;
  assign \new_Sorter100|15323_  = \new_Sorter100|15223_  & \new_Sorter100|15224_ ;
  assign \new_Sorter100|15324_  = \new_Sorter100|15223_  | \new_Sorter100|15224_ ;
  assign \new_Sorter100|15325_  = \new_Sorter100|15225_  & \new_Sorter100|15226_ ;
  assign \new_Sorter100|15326_  = \new_Sorter100|15225_  | \new_Sorter100|15226_ ;
  assign \new_Sorter100|15327_  = \new_Sorter100|15227_  & \new_Sorter100|15228_ ;
  assign \new_Sorter100|15328_  = \new_Sorter100|15227_  | \new_Sorter100|15228_ ;
  assign \new_Sorter100|15329_  = \new_Sorter100|15229_  & \new_Sorter100|15230_ ;
  assign \new_Sorter100|15330_  = \new_Sorter100|15229_  | \new_Sorter100|15230_ ;
  assign \new_Sorter100|15331_  = \new_Sorter100|15231_  & \new_Sorter100|15232_ ;
  assign \new_Sorter100|15332_  = \new_Sorter100|15231_  | \new_Sorter100|15232_ ;
  assign \new_Sorter100|15333_  = \new_Sorter100|15233_  & \new_Sorter100|15234_ ;
  assign \new_Sorter100|15334_  = \new_Sorter100|15233_  | \new_Sorter100|15234_ ;
  assign \new_Sorter100|15335_  = \new_Sorter100|15235_  & \new_Sorter100|15236_ ;
  assign \new_Sorter100|15336_  = \new_Sorter100|15235_  | \new_Sorter100|15236_ ;
  assign \new_Sorter100|15337_  = \new_Sorter100|15237_  & \new_Sorter100|15238_ ;
  assign \new_Sorter100|15338_  = \new_Sorter100|15237_  | \new_Sorter100|15238_ ;
  assign \new_Sorter100|15339_  = \new_Sorter100|15239_  & \new_Sorter100|15240_ ;
  assign \new_Sorter100|15340_  = \new_Sorter100|15239_  | \new_Sorter100|15240_ ;
  assign \new_Sorter100|15341_  = \new_Sorter100|15241_  & \new_Sorter100|15242_ ;
  assign \new_Sorter100|15342_  = \new_Sorter100|15241_  | \new_Sorter100|15242_ ;
  assign \new_Sorter100|15343_  = \new_Sorter100|15243_  & \new_Sorter100|15244_ ;
  assign \new_Sorter100|15344_  = \new_Sorter100|15243_  | \new_Sorter100|15244_ ;
  assign \new_Sorter100|15345_  = \new_Sorter100|15245_  & \new_Sorter100|15246_ ;
  assign \new_Sorter100|15346_  = \new_Sorter100|15245_  | \new_Sorter100|15246_ ;
  assign \new_Sorter100|15347_  = \new_Sorter100|15247_  & \new_Sorter100|15248_ ;
  assign \new_Sorter100|15348_  = \new_Sorter100|15247_  | \new_Sorter100|15248_ ;
  assign \new_Sorter100|15349_  = \new_Sorter100|15249_  & \new_Sorter100|15250_ ;
  assign \new_Sorter100|15350_  = \new_Sorter100|15249_  | \new_Sorter100|15250_ ;
  assign \new_Sorter100|15351_  = \new_Sorter100|15251_  & \new_Sorter100|15252_ ;
  assign \new_Sorter100|15352_  = \new_Sorter100|15251_  | \new_Sorter100|15252_ ;
  assign \new_Sorter100|15353_  = \new_Sorter100|15253_  & \new_Sorter100|15254_ ;
  assign \new_Sorter100|15354_  = \new_Sorter100|15253_  | \new_Sorter100|15254_ ;
  assign \new_Sorter100|15355_  = \new_Sorter100|15255_  & \new_Sorter100|15256_ ;
  assign \new_Sorter100|15356_  = \new_Sorter100|15255_  | \new_Sorter100|15256_ ;
  assign \new_Sorter100|15357_  = \new_Sorter100|15257_  & \new_Sorter100|15258_ ;
  assign \new_Sorter100|15358_  = \new_Sorter100|15257_  | \new_Sorter100|15258_ ;
  assign \new_Sorter100|15359_  = \new_Sorter100|15259_  & \new_Sorter100|15260_ ;
  assign \new_Sorter100|15360_  = \new_Sorter100|15259_  | \new_Sorter100|15260_ ;
  assign \new_Sorter100|15361_  = \new_Sorter100|15261_  & \new_Sorter100|15262_ ;
  assign \new_Sorter100|15362_  = \new_Sorter100|15261_  | \new_Sorter100|15262_ ;
  assign \new_Sorter100|15363_  = \new_Sorter100|15263_  & \new_Sorter100|15264_ ;
  assign \new_Sorter100|15364_  = \new_Sorter100|15263_  | \new_Sorter100|15264_ ;
  assign \new_Sorter100|15365_  = \new_Sorter100|15265_  & \new_Sorter100|15266_ ;
  assign \new_Sorter100|15366_  = \new_Sorter100|15265_  | \new_Sorter100|15266_ ;
  assign \new_Sorter100|15367_  = \new_Sorter100|15267_  & \new_Sorter100|15268_ ;
  assign \new_Sorter100|15368_  = \new_Sorter100|15267_  | \new_Sorter100|15268_ ;
  assign \new_Sorter100|15369_  = \new_Sorter100|15269_  & \new_Sorter100|15270_ ;
  assign \new_Sorter100|15370_  = \new_Sorter100|15269_  | \new_Sorter100|15270_ ;
  assign \new_Sorter100|15371_  = \new_Sorter100|15271_  & \new_Sorter100|15272_ ;
  assign \new_Sorter100|15372_  = \new_Sorter100|15271_  | \new_Sorter100|15272_ ;
  assign \new_Sorter100|15373_  = \new_Sorter100|15273_  & \new_Sorter100|15274_ ;
  assign \new_Sorter100|15374_  = \new_Sorter100|15273_  | \new_Sorter100|15274_ ;
  assign \new_Sorter100|15375_  = \new_Sorter100|15275_  & \new_Sorter100|15276_ ;
  assign \new_Sorter100|15376_  = \new_Sorter100|15275_  | \new_Sorter100|15276_ ;
  assign \new_Sorter100|15377_  = \new_Sorter100|15277_  & \new_Sorter100|15278_ ;
  assign \new_Sorter100|15378_  = \new_Sorter100|15277_  | \new_Sorter100|15278_ ;
  assign \new_Sorter100|15379_  = \new_Sorter100|15279_  & \new_Sorter100|15280_ ;
  assign \new_Sorter100|15380_  = \new_Sorter100|15279_  | \new_Sorter100|15280_ ;
  assign \new_Sorter100|15381_  = \new_Sorter100|15281_  & \new_Sorter100|15282_ ;
  assign \new_Sorter100|15382_  = \new_Sorter100|15281_  | \new_Sorter100|15282_ ;
  assign \new_Sorter100|15383_  = \new_Sorter100|15283_  & \new_Sorter100|15284_ ;
  assign \new_Sorter100|15384_  = \new_Sorter100|15283_  | \new_Sorter100|15284_ ;
  assign \new_Sorter100|15385_  = \new_Sorter100|15285_  & \new_Sorter100|15286_ ;
  assign \new_Sorter100|15386_  = \new_Sorter100|15285_  | \new_Sorter100|15286_ ;
  assign \new_Sorter100|15387_  = \new_Sorter100|15287_  & \new_Sorter100|15288_ ;
  assign \new_Sorter100|15388_  = \new_Sorter100|15287_  | \new_Sorter100|15288_ ;
  assign \new_Sorter100|15389_  = \new_Sorter100|15289_  & \new_Sorter100|15290_ ;
  assign \new_Sorter100|15390_  = \new_Sorter100|15289_  | \new_Sorter100|15290_ ;
  assign \new_Sorter100|15391_  = \new_Sorter100|15291_  & \new_Sorter100|15292_ ;
  assign \new_Sorter100|15392_  = \new_Sorter100|15291_  | \new_Sorter100|15292_ ;
  assign \new_Sorter100|15393_  = \new_Sorter100|15293_  & \new_Sorter100|15294_ ;
  assign \new_Sorter100|15394_  = \new_Sorter100|15293_  | \new_Sorter100|15294_ ;
  assign \new_Sorter100|15395_  = \new_Sorter100|15295_  & \new_Sorter100|15296_ ;
  assign \new_Sorter100|15396_  = \new_Sorter100|15295_  | \new_Sorter100|15296_ ;
  assign \new_Sorter100|15397_  = \new_Sorter100|15297_  & \new_Sorter100|15298_ ;
  assign \new_Sorter100|15398_  = \new_Sorter100|15297_  | \new_Sorter100|15298_ ;
  assign \new_Sorter100|15400_  = \new_Sorter100|15300_  & \new_Sorter100|15301_ ;
  assign \new_Sorter100|15401_  = \new_Sorter100|15300_  | \new_Sorter100|15301_ ;
  assign \new_Sorter100|15402_  = \new_Sorter100|15302_  & \new_Sorter100|15303_ ;
  assign \new_Sorter100|15403_  = \new_Sorter100|15302_  | \new_Sorter100|15303_ ;
  assign \new_Sorter100|15404_  = \new_Sorter100|15304_  & \new_Sorter100|15305_ ;
  assign \new_Sorter100|15405_  = \new_Sorter100|15304_  | \new_Sorter100|15305_ ;
  assign \new_Sorter100|15406_  = \new_Sorter100|15306_  & \new_Sorter100|15307_ ;
  assign \new_Sorter100|15407_  = \new_Sorter100|15306_  | \new_Sorter100|15307_ ;
  assign \new_Sorter100|15408_  = \new_Sorter100|15308_  & \new_Sorter100|15309_ ;
  assign \new_Sorter100|15409_  = \new_Sorter100|15308_  | \new_Sorter100|15309_ ;
  assign \new_Sorter100|15410_  = \new_Sorter100|15310_  & \new_Sorter100|15311_ ;
  assign \new_Sorter100|15411_  = \new_Sorter100|15310_  | \new_Sorter100|15311_ ;
  assign \new_Sorter100|15412_  = \new_Sorter100|15312_  & \new_Sorter100|15313_ ;
  assign \new_Sorter100|15413_  = \new_Sorter100|15312_  | \new_Sorter100|15313_ ;
  assign \new_Sorter100|15414_  = \new_Sorter100|15314_  & \new_Sorter100|15315_ ;
  assign \new_Sorter100|15415_  = \new_Sorter100|15314_  | \new_Sorter100|15315_ ;
  assign \new_Sorter100|15416_  = \new_Sorter100|15316_  & \new_Sorter100|15317_ ;
  assign \new_Sorter100|15417_  = \new_Sorter100|15316_  | \new_Sorter100|15317_ ;
  assign \new_Sorter100|15418_  = \new_Sorter100|15318_  & \new_Sorter100|15319_ ;
  assign \new_Sorter100|15419_  = \new_Sorter100|15318_  | \new_Sorter100|15319_ ;
  assign \new_Sorter100|15420_  = \new_Sorter100|15320_  & \new_Sorter100|15321_ ;
  assign \new_Sorter100|15421_  = \new_Sorter100|15320_  | \new_Sorter100|15321_ ;
  assign \new_Sorter100|15422_  = \new_Sorter100|15322_  & \new_Sorter100|15323_ ;
  assign \new_Sorter100|15423_  = \new_Sorter100|15322_  | \new_Sorter100|15323_ ;
  assign \new_Sorter100|15424_  = \new_Sorter100|15324_  & \new_Sorter100|15325_ ;
  assign \new_Sorter100|15425_  = \new_Sorter100|15324_  | \new_Sorter100|15325_ ;
  assign \new_Sorter100|15426_  = \new_Sorter100|15326_  & \new_Sorter100|15327_ ;
  assign \new_Sorter100|15427_  = \new_Sorter100|15326_  | \new_Sorter100|15327_ ;
  assign \new_Sorter100|15428_  = \new_Sorter100|15328_  & \new_Sorter100|15329_ ;
  assign \new_Sorter100|15429_  = \new_Sorter100|15328_  | \new_Sorter100|15329_ ;
  assign \new_Sorter100|15430_  = \new_Sorter100|15330_  & \new_Sorter100|15331_ ;
  assign \new_Sorter100|15431_  = \new_Sorter100|15330_  | \new_Sorter100|15331_ ;
  assign \new_Sorter100|15432_  = \new_Sorter100|15332_  & \new_Sorter100|15333_ ;
  assign \new_Sorter100|15433_  = \new_Sorter100|15332_  | \new_Sorter100|15333_ ;
  assign \new_Sorter100|15434_  = \new_Sorter100|15334_  & \new_Sorter100|15335_ ;
  assign \new_Sorter100|15435_  = \new_Sorter100|15334_  | \new_Sorter100|15335_ ;
  assign \new_Sorter100|15436_  = \new_Sorter100|15336_  & \new_Sorter100|15337_ ;
  assign \new_Sorter100|15437_  = \new_Sorter100|15336_  | \new_Sorter100|15337_ ;
  assign \new_Sorter100|15438_  = \new_Sorter100|15338_  & \new_Sorter100|15339_ ;
  assign \new_Sorter100|15439_  = \new_Sorter100|15338_  | \new_Sorter100|15339_ ;
  assign \new_Sorter100|15440_  = \new_Sorter100|15340_  & \new_Sorter100|15341_ ;
  assign \new_Sorter100|15441_  = \new_Sorter100|15340_  | \new_Sorter100|15341_ ;
  assign \new_Sorter100|15442_  = \new_Sorter100|15342_  & \new_Sorter100|15343_ ;
  assign \new_Sorter100|15443_  = \new_Sorter100|15342_  | \new_Sorter100|15343_ ;
  assign \new_Sorter100|15444_  = \new_Sorter100|15344_  & \new_Sorter100|15345_ ;
  assign \new_Sorter100|15445_  = \new_Sorter100|15344_  | \new_Sorter100|15345_ ;
  assign \new_Sorter100|15446_  = \new_Sorter100|15346_  & \new_Sorter100|15347_ ;
  assign \new_Sorter100|15447_  = \new_Sorter100|15346_  | \new_Sorter100|15347_ ;
  assign \new_Sorter100|15448_  = \new_Sorter100|15348_  & \new_Sorter100|15349_ ;
  assign \new_Sorter100|15449_  = \new_Sorter100|15348_  | \new_Sorter100|15349_ ;
  assign \new_Sorter100|15450_  = \new_Sorter100|15350_  & \new_Sorter100|15351_ ;
  assign \new_Sorter100|15451_  = \new_Sorter100|15350_  | \new_Sorter100|15351_ ;
  assign \new_Sorter100|15452_  = \new_Sorter100|15352_  & \new_Sorter100|15353_ ;
  assign \new_Sorter100|15453_  = \new_Sorter100|15352_  | \new_Sorter100|15353_ ;
  assign \new_Sorter100|15454_  = \new_Sorter100|15354_  & \new_Sorter100|15355_ ;
  assign \new_Sorter100|15455_  = \new_Sorter100|15354_  | \new_Sorter100|15355_ ;
  assign \new_Sorter100|15456_  = \new_Sorter100|15356_  & \new_Sorter100|15357_ ;
  assign \new_Sorter100|15457_  = \new_Sorter100|15356_  | \new_Sorter100|15357_ ;
  assign \new_Sorter100|15458_  = \new_Sorter100|15358_  & \new_Sorter100|15359_ ;
  assign \new_Sorter100|15459_  = \new_Sorter100|15358_  | \new_Sorter100|15359_ ;
  assign \new_Sorter100|15460_  = \new_Sorter100|15360_  & \new_Sorter100|15361_ ;
  assign \new_Sorter100|15461_  = \new_Sorter100|15360_  | \new_Sorter100|15361_ ;
  assign \new_Sorter100|15462_  = \new_Sorter100|15362_  & \new_Sorter100|15363_ ;
  assign \new_Sorter100|15463_  = \new_Sorter100|15362_  | \new_Sorter100|15363_ ;
  assign \new_Sorter100|15464_  = \new_Sorter100|15364_  & \new_Sorter100|15365_ ;
  assign \new_Sorter100|15465_  = \new_Sorter100|15364_  | \new_Sorter100|15365_ ;
  assign \new_Sorter100|15466_  = \new_Sorter100|15366_  & \new_Sorter100|15367_ ;
  assign \new_Sorter100|15467_  = \new_Sorter100|15366_  | \new_Sorter100|15367_ ;
  assign \new_Sorter100|15468_  = \new_Sorter100|15368_  & \new_Sorter100|15369_ ;
  assign \new_Sorter100|15469_  = \new_Sorter100|15368_  | \new_Sorter100|15369_ ;
  assign \new_Sorter100|15470_  = \new_Sorter100|15370_  & \new_Sorter100|15371_ ;
  assign \new_Sorter100|15471_  = \new_Sorter100|15370_  | \new_Sorter100|15371_ ;
  assign \new_Sorter100|15472_  = \new_Sorter100|15372_  & \new_Sorter100|15373_ ;
  assign \new_Sorter100|15473_  = \new_Sorter100|15372_  | \new_Sorter100|15373_ ;
  assign \new_Sorter100|15474_  = \new_Sorter100|15374_  & \new_Sorter100|15375_ ;
  assign \new_Sorter100|15475_  = \new_Sorter100|15374_  | \new_Sorter100|15375_ ;
  assign \new_Sorter100|15476_  = \new_Sorter100|15376_  & \new_Sorter100|15377_ ;
  assign \new_Sorter100|15477_  = \new_Sorter100|15376_  | \new_Sorter100|15377_ ;
  assign \new_Sorter100|15478_  = \new_Sorter100|15378_  & \new_Sorter100|15379_ ;
  assign \new_Sorter100|15479_  = \new_Sorter100|15378_  | \new_Sorter100|15379_ ;
  assign \new_Sorter100|15480_  = \new_Sorter100|15380_  & \new_Sorter100|15381_ ;
  assign \new_Sorter100|15481_  = \new_Sorter100|15380_  | \new_Sorter100|15381_ ;
  assign \new_Sorter100|15482_  = \new_Sorter100|15382_  & \new_Sorter100|15383_ ;
  assign \new_Sorter100|15483_  = \new_Sorter100|15382_  | \new_Sorter100|15383_ ;
  assign \new_Sorter100|15484_  = \new_Sorter100|15384_  & \new_Sorter100|15385_ ;
  assign \new_Sorter100|15485_  = \new_Sorter100|15384_  | \new_Sorter100|15385_ ;
  assign \new_Sorter100|15486_  = \new_Sorter100|15386_  & \new_Sorter100|15387_ ;
  assign \new_Sorter100|15487_  = \new_Sorter100|15386_  | \new_Sorter100|15387_ ;
  assign \new_Sorter100|15488_  = \new_Sorter100|15388_  & \new_Sorter100|15389_ ;
  assign \new_Sorter100|15489_  = \new_Sorter100|15388_  | \new_Sorter100|15389_ ;
  assign \new_Sorter100|15490_  = \new_Sorter100|15390_  & \new_Sorter100|15391_ ;
  assign \new_Sorter100|15491_  = \new_Sorter100|15390_  | \new_Sorter100|15391_ ;
  assign \new_Sorter100|15492_  = \new_Sorter100|15392_  & \new_Sorter100|15393_ ;
  assign \new_Sorter100|15493_  = \new_Sorter100|15392_  | \new_Sorter100|15393_ ;
  assign \new_Sorter100|15494_  = \new_Sorter100|15394_  & \new_Sorter100|15395_ ;
  assign \new_Sorter100|15495_  = \new_Sorter100|15394_  | \new_Sorter100|15395_ ;
  assign \new_Sorter100|15496_  = \new_Sorter100|15396_  & \new_Sorter100|15397_ ;
  assign \new_Sorter100|15497_  = \new_Sorter100|15396_  | \new_Sorter100|15397_ ;
  assign \new_Sorter100|15498_  = \new_Sorter100|15398_  & \new_Sorter100|15399_ ;
  assign \new_Sorter100|15499_  = \new_Sorter100|15398_  | \new_Sorter100|15399_ ;
  assign \new_Sorter100|15500_  = \new_Sorter100|15400_ ;
  assign \new_Sorter100|15599_  = \new_Sorter100|15499_ ;
  assign \new_Sorter100|15501_  = \new_Sorter100|15401_  & \new_Sorter100|15402_ ;
  assign \new_Sorter100|15502_  = \new_Sorter100|15401_  | \new_Sorter100|15402_ ;
  assign \new_Sorter100|15503_  = \new_Sorter100|15403_  & \new_Sorter100|15404_ ;
  assign \new_Sorter100|15504_  = \new_Sorter100|15403_  | \new_Sorter100|15404_ ;
  assign \new_Sorter100|15505_  = \new_Sorter100|15405_  & \new_Sorter100|15406_ ;
  assign \new_Sorter100|15506_  = \new_Sorter100|15405_  | \new_Sorter100|15406_ ;
  assign \new_Sorter100|15507_  = \new_Sorter100|15407_  & \new_Sorter100|15408_ ;
  assign \new_Sorter100|15508_  = \new_Sorter100|15407_  | \new_Sorter100|15408_ ;
  assign \new_Sorter100|15509_  = \new_Sorter100|15409_  & \new_Sorter100|15410_ ;
  assign \new_Sorter100|15510_  = \new_Sorter100|15409_  | \new_Sorter100|15410_ ;
  assign \new_Sorter100|15511_  = \new_Sorter100|15411_  & \new_Sorter100|15412_ ;
  assign \new_Sorter100|15512_  = \new_Sorter100|15411_  | \new_Sorter100|15412_ ;
  assign \new_Sorter100|15513_  = \new_Sorter100|15413_  & \new_Sorter100|15414_ ;
  assign \new_Sorter100|15514_  = \new_Sorter100|15413_  | \new_Sorter100|15414_ ;
  assign \new_Sorter100|15515_  = \new_Sorter100|15415_  & \new_Sorter100|15416_ ;
  assign \new_Sorter100|15516_  = \new_Sorter100|15415_  | \new_Sorter100|15416_ ;
  assign \new_Sorter100|15517_  = \new_Sorter100|15417_  & \new_Sorter100|15418_ ;
  assign \new_Sorter100|15518_  = \new_Sorter100|15417_  | \new_Sorter100|15418_ ;
  assign \new_Sorter100|15519_  = \new_Sorter100|15419_  & \new_Sorter100|15420_ ;
  assign \new_Sorter100|15520_  = \new_Sorter100|15419_  | \new_Sorter100|15420_ ;
  assign \new_Sorter100|15521_  = \new_Sorter100|15421_  & \new_Sorter100|15422_ ;
  assign \new_Sorter100|15522_  = \new_Sorter100|15421_  | \new_Sorter100|15422_ ;
  assign \new_Sorter100|15523_  = \new_Sorter100|15423_  & \new_Sorter100|15424_ ;
  assign \new_Sorter100|15524_  = \new_Sorter100|15423_  | \new_Sorter100|15424_ ;
  assign \new_Sorter100|15525_  = \new_Sorter100|15425_  & \new_Sorter100|15426_ ;
  assign \new_Sorter100|15526_  = \new_Sorter100|15425_  | \new_Sorter100|15426_ ;
  assign \new_Sorter100|15527_  = \new_Sorter100|15427_  & \new_Sorter100|15428_ ;
  assign \new_Sorter100|15528_  = \new_Sorter100|15427_  | \new_Sorter100|15428_ ;
  assign \new_Sorter100|15529_  = \new_Sorter100|15429_  & \new_Sorter100|15430_ ;
  assign \new_Sorter100|15530_  = \new_Sorter100|15429_  | \new_Sorter100|15430_ ;
  assign \new_Sorter100|15531_  = \new_Sorter100|15431_  & \new_Sorter100|15432_ ;
  assign \new_Sorter100|15532_  = \new_Sorter100|15431_  | \new_Sorter100|15432_ ;
  assign \new_Sorter100|15533_  = \new_Sorter100|15433_  & \new_Sorter100|15434_ ;
  assign \new_Sorter100|15534_  = \new_Sorter100|15433_  | \new_Sorter100|15434_ ;
  assign \new_Sorter100|15535_  = \new_Sorter100|15435_  & \new_Sorter100|15436_ ;
  assign \new_Sorter100|15536_  = \new_Sorter100|15435_  | \new_Sorter100|15436_ ;
  assign \new_Sorter100|15537_  = \new_Sorter100|15437_  & \new_Sorter100|15438_ ;
  assign \new_Sorter100|15538_  = \new_Sorter100|15437_  | \new_Sorter100|15438_ ;
  assign \new_Sorter100|15539_  = \new_Sorter100|15439_  & \new_Sorter100|15440_ ;
  assign \new_Sorter100|15540_  = \new_Sorter100|15439_  | \new_Sorter100|15440_ ;
  assign \new_Sorter100|15541_  = \new_Sorter100|15441_  & \new_Sorter100|15442_ ;
  assign \new_Sorter100|15542_  = \new_Sorter100|15441_  | \new_Sorter100|15442_ ;
  assign \new_Sorter100|15543_  = \new_Sorter100|15443_  & \new_Sorter100|15444_ ;
  assign \new_Sorter100|15544_  = \new_Sorter100|15443_  | \new_Sorter100|15444_ ;
  assign \new_Sorter100|15545_  = \new_Sorter100|15445_  & \new_Sorter100|15446_ ;
  assign \new_Sorter100|15546_  = \new_Sorter100|15445_  | \new_Sorter100|15446_ ;
  assign \new_Sorter100|15547_  = \new_Sorter100|15447_  & \new_Sorter100|15448_ ;
  assign \new_Sorter100|15548_  = \new_Sorter100|15447_  | \new_Sorter100|15448_ ;
  assign \new_Sorter100|15549_  = \new_Sorter100|15449_  & \new_Sorter100|15450_ ;
  assign \new_Sorter100|15550_  = \new_Sorter100|15449_  | \new_Sorter100|15450_ ;
  assign \new_Sorter100|15551_  = \new_Sorter100|15451_  & \new_Sorter100|15452_ ;
  assign \new_Sorter100|15552_  = \new_Sorter100|15451_  | \new_Sorter100|15452_ ;
  assign \new_Sorter100|15553_  = \new_Sorter100|15453_  & \new_Sorter100|15454_ ;
  assign \new_Sorter100|15554_  = \new_Sorter100|15453_  | \new_Sorter100|15454_ ;
  assign \new_Sorter100|15555_  = \new_Sorter100|15455_  & \new_Sorter100|15456_ ;
  assign \new_Sorter100|15556_  = \new_Sorter100|15455_  | \new_Sorter100|15456_ ;
  assign \new_Sorter100|15557_  = \new_Sorter100|15457_  & \new_Sorter100|15458_ ;
  assign \new_Sorter100|15558_  = \new_Sorter100|15457_  | \new_Sorter100|15458_ ;
  assign \new_Sorter100|15559_  = \new_Sorter100|15459_  & \new_Sorter100|15460_ ;
  assign \new_Sorter100|15560_  = \new_Sorter100|15459_  | \new_Sorter100|15460_ ;
  assign \new_Sorter100|15561_  = \new_Sorter100|15461_  & \new_Sorter100|15462_ ;
  assign \new_Sorter100|15562_  = \new_Sorter100|15461_  | \new_Sorter100|15462_ ;
  assign \new_Sorter100|15563_  = \new_Sorter100|15463_  & \new_Sorter100|15464_ ;
  assign \new_Sorter100|15564_  = \new_Sorter100|15463_  | \new_Sorter100|15464_ ;
  assign \new_Sorter100|15565_  = \new_Sorter100|15465_  & \new_Sorter100|15466_ ;
  assign \new_Sorter100|15566_  = \new_Sorter100|15465_  | \new_Sorter100|15466_ ;
  assign \new_Sorter100|15567_  = \new_Sorter100|15467_  & \new_Sorter100|15468_ ;
  assign \new_Sorter100|15568_  = \new_Sorter100|15467_  | \new_Sorter100|15468_ ;
  assign \new_Sorter100|15569_  = \new_Sorter100|15469_  & \new_Sorter100|15470_ ;
  assign \new_Sorter100|15570_  = \new_Sorter100|15469_  | \new_Sorter100|15470_ ;
  assign \new_Sorter100|15571_  = \new_Sorter100|15471_  & \new_Sorter100|15472_ ;
  assign \new_Sorter100|15572_  = \new_Sorter100|15471_  | \new_Sorter100|15472_ ;
  assign \new_Sorter100|15573_  = \new_Sorter100|15473_  & \new_Sorter100|15474_ ;
  assign \new_Sorter100|15574_  = \new_Sorter100|15473_  | \new_Sorter100|15474_ ;
  assign \new_Sorter100|15575_  = \new_Sorter100|15475_  & \new_Sorter100|15476_ ;
  assign \new_Sorter100|15576_  = \new_Sorter100|15475_  | \new_Sorter100|15476_ ;
  assign \new_Sorter100|15577_  = \new_Sorter100|15477_  & \new_Sorter100|15478_ ;
  assign \new_Sorter100|15578_  = \new_Sorter100|15477_  | \new_Sorter100|15478_ ;
  assign \new_Sorter100|15579_  = \new_Sorter100|15479_  & \new_Sorter100|15480_ ;
  assign \new_Sorter100|15580_  = \new_Sorter100|15479_  | \new_Sorter100|15480_ ;
  assign \new_Sorter100|15581_  = \new_Sorter100|15481_  & \new_Sorter100|15482_ ;
  assign \new_Sorter100|15582_  = \new_Sorter100|15481_  | \new_Sorter100|15482_ ;
  assign \new_Sorter100|15583_  = \new_Sorter100|15483_  & \new_Sorter100|15484_ ;
  assign \new_Sorter100|15584_  = \new_Sorter100|15483_  | \new_Sorter100|15484_ ;
  assign \new_Sorter100|15585_  = \new_Sorter100|15485_  & \new_Sorter100|15486_ ;
  assign \new_Sorter100|15586_  = \new_Sorter100|15485_  | \new_Sorter100|15486_ ;
  assign \new_Sorter100|15587_  = \new_Sorter100|15487_  & \new_Sorter100|15488_ ;
  assign \new_Sorter100|15588_  = \new_Sorter100|15487_  | \new_Sorter100|15488_ ;
  assign \new_Sorter100|15589_  = \new_Sorter100|15489_  & \new_Sorter100|15490_ ;
  assign \new_Sorter100|15590_  = \new_Sorter100|15489_  | \new_Sorter100|15490_ ;
  assign \new_Sorter100|15591_  = \new_Sorter100|15491_  & \new_Sorter100|15492_ ;
  assign \new_Sorter100|15592_  = \new_Sorter100|15491_  | \new_Sorter100|15492_ ;
  assign \new_Sorter100|15593_  = \new_Sorter100|15493_  & \new_Sorter100|15494_ ;
  assign \new_Sorter100|15594_  = \new_Sorter100|15493_  | \new_Sorter100|15494_ ;
  assign \new_Sorter100|15595_  = \new_Sorter100|15495_  & \new_Sorter100|15496_ ;
  assign \new_Sorter100|15596_  = \new_Sorter100|15495_  | \new_Sorter100|15496_ ;
  assign \new_Sorter100|15597_  = \new_Sorter100|15497_  & \new_Sorter100|15498_ ;
  assign \new_Sorter100|15598_  = \new_Sorter100|15497_  | \new_Sorter100|15498_ ;
  assign \new_Sorter100|15600_  = \new_Sorter100|15500_  & \new_Sorter100|15501_ ;
  assign \new_Sorter100|15601_  = \new_Sorter100|15500_  | \new_Sorter100|15501_ ;
  assign \new_Sorter100|15602_  = \new_Sorter100|15502_  & \new_Sorter100|15503_ ;
  assign \new_Sorter100|15603_  = \new_Sorter100|15502_  | \new_Sorter100|15503_ ;
  assign \new_Sorter100|15604_  = \new_Sorter100|15504_  & \new_Sorter100|15505_ ;
  assign \new_Sorter100|15605_  = \new_Sorter100|15504_  | \new_Sorter100|15505_ ;
  assign \new_Sorter100|15606_  = \new_Sorter100|15506_  & \new_Sorter100|15507_ ;
  assign \new_Sorter100|15607_  = \new_Sorter100|15506_  | \new_Sorter100|15507_ ;
  assign \new_Sorter100|15608_  = \new_Sorter100|15508_  & \new_Sorter100|15509_ ;
  assign \new_Sorter100|15609_  = \new_Sorter100|15508_  | \new_Sorter100|15509_ ;
  assign \new_Sorter100|15610_  = \new_Sorter100|15510_  & \new_Sorter100|15511_ ;
  assign \new_Sorter100|15611_  = \new_Sorter100|15510_  | \new_Sorter100|15511_ ;
  assign \new_Sorter100|15612_  = \new_Sorter100|15512_  & \new_Sorter100|15513_ ;
  assign \new_Sorter100|15613_  = \new_Sorter100|15512_  | \new_Sorter100|15513_ ;
  assign \new_Sorter100|15614_  = \new_Sorter100|15514_  & \new_Sorter100|15515_ ;
  assign \new_Sorter100|15615_  = \new_Sorter100|15514_  | \new_Sorter100|15515_ ;
  assign \new_Sorter100|15616_  = \new_Sorter100|15516_  & \new_Sorter100|15517_ ;
  assign \new_Sorter100|15617_  = \new_Sorter100|15516_  | \new_Sorter100|15517_ ;
  assign \new_Sorter100|15618_  = \new_Sorter100|15518_  & \new_Sorter100|15519_ ;
  assign \new_Sorter100|15619_  = \new_Sorter100|15518_  | \new_Sorter100|15519_ ;
  assign \new_Sorter100|15620_  = \new_Sorter100|15520_  & \new_Sorter100|15521_ ;
  assign \new_Sorter100|15621_  = \new_Sorter100|15520_  | \new_Sorter100|15521_ ;
  assign \new_Sorter100|15622_  = \new_Sorter100|15522_  & \new_Sorter100|15523_ ;
  assign \new_Sorter100|15623_  = \new_Sorter100|15522_  | \new_Sorter100|15523_ ;
  assign \new_Sorter100|15624_  = \new_Sorter100|15524_  & \new_Sorter100|15525_ ;
  assign \new_Sorter100|15625_  = \new_Sorter100|15524_  | \new_Sorter100|15525_ ;
  assign \new_Sorter100|15626_  = \new_Sorter100|15526_  & \new_Sorter100|15527_ ;
  assign \new_Sorter100|15627_  = \new_Sorter100|15526_  | \new_Sorter100|15527_ ;
  assign \new_Sorter100|15628_  = \new_Sorter100|15528_  & \new_Sorter100|15529_ ;
  assign \new_Sorter100|15629_  = \new_Sorter100|15528_  | \new_Sorter100|15529_ ;
  assign \new_Sorter100|15630_  = \new_Sorter100|15530_  & \new_Sorter100|15531_ ;
  assign \new_Sorter100|15631_  = \new_Sorter100|15530_  | \new_Sorter100|15531_ ;
  assign \new_Sorter100|15632_  = \new_Sorter100|15532_  & \new_Sorter100|15533_ ;
  assign \new_Sorter100|15633_  = \new_Sorter100|15532_  | \new_Sorter100|15533_ ;
  assign \new_Sorter100|15634_  = \new_Sorter100|15534_  & \new_Sorter100|15535_ ;
  assign \new_Sorter100|15635_  = \new_Sorter100|15534_  | \new_Sorter100|15535_ ;
  assign \new_Sorter100|15636_  = \new_Sorter100|15536_  & \new_Sorter100|15537_ ;
  assign \new_Sorter100|15637_  = \new_Sorter100|15536_  | \new_Sorter100|15537_ ;
  assign \new_Sorter100|15638_  = \new_Sorter100|15538_  & \new_Sorter100|15539_ ;
  assign \new_Sorter100|15639_  = \new_Sorter100|15538_  | \new_Sorter100|15539_ ;
  assign \new_Sorter100|15640_  = \new_Sorter100|15540_  & \new_Sorter100|15541_ ;
  assign \new_Sorter100|15641_  = \new_Sorter100|15540_  | \new_Sorter100|15541_ ;
  assign \new_Sorter100|15642_  = \new_Sorter100|15542_  & \new_Sorter100|15543_ ;
  assign \new_Sorter100|15643_  = \new_Sorter100|15542_  | \new_Sorter100|15543_ ;
  assign \new_Sorter100|15644_  = \new_Sorter100|15544_  & \new_Sorter100|15545_ ;
  assign \new_Sorter100|15645_  = \new_Sorter100|15544_  | \new_Sorter100|15545_ ;
  assign \new_Sorter100|15646_  = \new_Sorter100|15546_  & \new_Sorter100|15547_ ;
  assign \new_Sorter100|15647_  = \new_Sorter100|15546_  | \new_Sorter100|15547_ ;
  assign \new_Sorter100|15648_  = \new_Sorter100|15548_  & \new_Sorter100|15549_ ;
  assign \new_Sorter100|15649_  = \new_Sorter100|15548_  | \new_Sorter100|15549_ ;
  assign \new_Sorter100|15650_  = \new_Sorter100|15550_  & \new_Sorter100|15551_ ;
  assign \new_Sorter100|15651_  = \new_Sorter100|15550_  | \new_Sorter100|15551_ ;
  assign \new_Sorter100|15652_  = \new_Sorter100|15552_  & \new_Sorter100|15553_ ;
  assign \new_Sorter100|15653_  = \new_Sorter100|15552_  | \new_Sorter100|15553_ ;
  assign \new_Sorter100|15654_  = \new_Sorter100|15554_  & \new_Sorter100|15555_ ;
  assign \new_Sorter100|15655_  = \new_Sorter100|15554_  | \new_Sorter100|15555_ ;
  assign \new_Sorter100|15656_  = \new_Sorter100|15556_  & \new_Sorter100|15557_ ;
  assign \new_Sorter100|15657_  = \new_Sorter100|15556_  | \new_Sorter100|15557_ ;
  assign \new_Sorter100|15658_  = \new_Sorter100|15558_  & \new_Sorter100|15559_ ;
  assign \new_Sorter100|15659_  = \new_Sorter100|15558_  | \new_Sorter100|15559_ ;
  assign \new_Sorter100|15660_  = \new_Sorter100|15560_  & \new_Sorter100|15561_ ;
  assign \new_Sorter100|15661_  = \new_Sorter100|15560_  | \new_Sorter100|15561_ ;
  assign \new_Sorter100|15662_  = \new_Sorter100|15562_  & \new_Sorter100|15563_ ;
  assign \new_Sorter100|15663_  = \new_Sorter100|15562_  | \new_Sorter100|15563_ ;
  assign \new_Sorter100|15664_  = \new_Sorter100|15564_  & \new_Sorter100|15565_ ;
  assign \new_Sorter100|15665_  = \new_Sorter100|15564_  | \new_Sorter100|15565_ ;
  assign \new_Sorter100|15666_  = \new_Sorter100|15566_  & \new_Sorter100|15567_ ;
  assign \new_Sorter100|15667_  = \new_Sorter100|15566_  | \new_Sorter100|15567_ ;
  assign \new_Sorter100|15668_  = \new_Sorter100|15568_  & \new_Sorter100|15569_ ;
  assign \new_Sorter100|15669_  = \new_Sorter100|15568_  | \new_Sorter100|15569_ ;
  assign \new_Sorter100|15670_  = \new_Sorter100|15570_  & \new_Sorter100|15571_ ;
  assign \new_Sorter100|15671_  = \new_Sorter100|15570_  | \new_Sorter100|15571_ ;
  assign \new_Sorter100|15672_  = \new_Sorter100|15572_  & \new_Sorter100|15573_ ;
  assign \new_Sorter100|15673_  = \new_Sorter100|15572_  | \new_Sorter100|15573_ ;
  assign \new_Sorter100|15674_  = \new_Sorter100|15574_  & \new_Sorter100|15575_ ;
  assign \new_Sorter100|15675_  = \new_Sorter100|15574_  | \new_Sorter100|15575_ ;
  assign \new_Sorter100|15676_  = \new_Sorter100|15576_  & \new_Sorter100|15577_ ;
  assign \new_Sorter100|15677_  = \new_Sorter100|15576_  | \new_Sorter100|15577_ ;
  assign \new_Sorter100|15678_  = \new_Sorter100|15578_  & \new_Sorter100|15579_ ;
  assign \new_Sorter100|15679_  = \new_Sorter100|15578_  | \new_Sorter100|15579_ ;
  assign \new_Sorter100|15680_  = \new_Sorter100|15580_  & \new_Sorter100|15581_ ;
  assign \new_Sorter100|15681_  = \new_Sorter100|15580_  | \new_Sorter100|15581_ ;
  assign \new_Sorter100|15682_  = \new_Sorter100|15582_  & \new_Sorter100|15583_ ;
  assign \new_Sorter100|15683_  = \new_Sorter100|15582_  | \new_Sorter100|15583_ ;
  assign \new_Sorter100|15684_  = \new_Sorter100|15584_  & \new_Sorter100|15585_ ;
  assign \new_Sorter100|15685_  = \new_Sorter100|15584_  | \new_Sorter100|15585_ ;
  assign \new_Sorter100|15686_  = \new_Sorter100|15586_  & \new_Sorter100|15587_ ;
  assign \new_Sorter100|15687_  = \new_Sorter100|15586_  | \new_Sorter100|15587_ ;
  assign \new_Sorter100|15688_  = \new_Sorter100|15588_  & \new_Sorter100|15589_ ;
  assign \new_Sorter100|15689_  = \new_Sorter100|15588_  | \new_Sorter100|15589_ ;
  assign \new_Sorter100|15690_  = \new_Sorter100|15590_  & \new_Sorter100|15591_ ;
  assign \new_Sorter100|15691_  = \new_Sorter100|15590_  | \new_Sorter100|15591_ ;
  assign \new_Sorter100|15692_  = \new_Sorter100|15592_  & \new_Sorter100|15593_ ;
  assign \new_Sorter100|15693_  = \new_Sorter100|15592_  | \new_Sorter100|15593_ ;
  assign \new_Sorter100|15694_  = \new_Sorter100|15594_  & \new_Sorter100|15595_ ;
  assign \new_Sorter100|15695_  = \new_Sorter100|15594_  | \new_Sorter100|15595_ ;
  assign \new_Sorter100|15696_  = \new_Sorter100|15596_  & \new_Sorter100|15597_ ;
  assign \new_Sorter100|15697_  = \new_Sorter100|15596_  | \new_Sorter100|15597_ ;
  assign \new_Sorter100|15698_  = \new_Sorter100|15598_  & \new_Sorter100|15599_ ;
  assign \new_Sorter100|15699_  = \new_Sorter100|15598_  | \new_Sorter100|15599_ ;
  assign \new_Sorter100|15700_  = \new_Sorter100|15600_ ;
  assign \new_Sorter100|15799_  = \new_Sorter100|15699_ ;
  assign \new_Sorter100|15701_  = \new_Sorter100|15601_  & \new_Sorter100|15602_ ;
  assign \new_Sorter100|15702_  = \new_Sorter100|15601_  | \new_Sorter100|15602_ ;
  assign \new_Sorter100|15703_  = \new_Sorter100|15603_  & \new_Sorter100|15604_ ;
  assign \new_Sorter100|15704_  = \new_Sorter100|15603_  | \new_Sorter100|15604_ ;
  assign \new_Sorter100|15705_  = \new_Sorter100|15605_  & \new_Sorter100|15606_ ;
  assign \new_Sorter100|15706_  = \new_Sorter100|15605_  | \new_Sorter100|15606_ ;
  assign \new_Sorter100|15707_  = \new_Sorter100|15607_  & \new_Sorter100|15608_ ;
  assign \new_Sorter100|15708_  = \new_Sorter100|15607_  | \new_Sorter100|15608_ ;
  assign \new_Sorter100|15709_  = \new_Sorter100|15609_  & \new_Sorter100|15610_ ;
  assign \new_Sorter100|15710_  = \new_Sorter100|15609_  | \new_Sorter100|15610_ ;
  assign \new_Sorter100|15711_  = \new_Sorter100|15611_  & \new_Sorter100|15612_ ;
  assign \new_Sorter100|15712_  = \new_Sorter100|15611_  | \new_Sorter100|15612_ ;
  assign \new_Sorter100|15713_  = \new_Sorter100|15613_  & \new_Sorter100|15614_ ;
  assign \new_Sorter100|15714_  = \new_Sorter100|15613_  | \new_Sorter100|15614_ ;
  assign \new_Sorter100|15715_  = \new_Sorter100|15615_  & \new_Sorter100|15616_ ;
  assign \new_Sorter100|15716_  = \new_Sorter100|15615_  | \new_Sorter100|15616_ ;
  assign \new_Sorter100|15717_  = \new_Sorter100|15617_  & \new_Sorter100|15618_ ;
  assign \new_Sorter100|15718_  = \new_Sorter100|15617_  | \new_Sorter100|15618_ ;
  assign \new_Sorter100|15719_  = \new_Sorter100|15619_  & \new_Sorter100|15620_ ;
  assign \new_Sorter100|15720_  = \new_Sorter100|15619_  | \new_Sorter100|15620_ ;
  assign \new_Sorter100|15721_  = \new_Sorter100|15621_  & \new_Sorter100|15622_ ;
  assign \new_Sorter100|15722_  = \new_Sorter100|15621_  | \new_Sorter100|15622_ ;
  assign \new_Sorter100|15723_  = \new_Sorter100|15623_  & \new_Sorter100|15624_ ;
  assign \new_Sorter100|15724_  = \new_Sorter100|15623_  | \new_Sorter100|15624_ ;
  assign \new_Sorter100|15725_  = \new_Sorter100|15625_  & \new_Sorter100|15626_ ;
  assign \new_Sorter100|15726_  = \new_Sorter100|15625_  | \new_Sorter100|15626_ ;
  assign \new_Sorter100|15727_  = \new_Sorter100|15627_  & \new_Sorter100|15628_ ;
  assign \new_Sorter100|15728_  = \new_Sorter100|15627_  | \new_Sorter100|15628_ ;
  assign \new_Sorter100|15729_  = \new_Sorter100|15629_  & \new_Sorter100|15630_ ;
  assign \new_Sorter100|15730_  = \new_Sorter100|15629_  | \new_Sorter100|15630_ ;
  assign \new_Sorter100|15731_  = \new_Sorter100|15631_  & \new_Sorter100|15632_ ;
  assign \new_Sorter100|15732_  = \new_Sorter100|15631_  | \new_Sorter100|15632_ ;
  assign \new_Sorter100|15733_  = \new_Sorter100|15633_  & \new_Sorter100|15634_ ;
  assign \new_Sorter100|15734_  = \new_Sorter100|15633_  | \new_Sorter100|15634_ ;
  assign \new_Sorter100|15735_  = \new_Sorter100|15635_  & \new_Sorter100|15636_ ;
  assign \new_Sorter100|15736_  = \new_Sorter100|15635_  | \new_Sorter100|15636_ ;
  assign \new_Sorter100|15737_  = \new_Sorter100|15637_  & \new_Sorter100|15638_ ;
  assign \new_Sorter100|15738_  = \new_Sorter100|15637_  | \new_Sorter100|15638_ ;
  assign \new_Sorter100|15739_  = \new_Sorter100|15639_  & \new_Sorter100|15640_ ;
  assign \new_Sorter100|15740_  = \new_Sorter100|15639_  | \new_Sorter100|15640_ ;
  assign \new_Sorter100|15741_  = \new_Sorter100|15641_  & \new_Sorter100|15642_ ;
  assign \new_Sorter100|15742_  = \new_Sorter100|15641_  | \new_Sorter100|15642_ ;
  assign \new_Sorter100|15743_  = \new_Sorter100|15643_  & \new_Sorter100|15644_ ;
  assign \new_Sorter100|15744_  = \new_Sorter100|15643_  | \new_Sorter100|15644_ ;
  assign \new_Sorter100|15745_  = \new_Sorter100|15645_  & \new_Sorter100|15646_ ;
  assign \new_Sorter100|15746_  = \new_Sorter100|15645_  | \new_Sorter100|15646_ ;
  assign \new_Sorter100|15747_  = \new_Sorter100|15647_  & \new_Sorter100|15648_ ;
  assign \new_Sorter100|15748_  = \new_Sorter100|15647_  | \new_Sorter100|15648_ ;
  assign \new_Sorter100|15749_  = \new_Sorter100|15649_  & \new_Sorter100|15650_ ;
  assign \new_Sorter100|15750_  = \new_Sorter100|15649_  | \new_Sorter100|15650_ ;
  assign \new_Sorter100|15751_  = \new_Sorter100|15651_  & \new_Sorter100|15652_ ;
  assign \new_Sorter100|15752_  = \new_Sorter100|15651_  | \new_Sorter100|15652_ ;
  assign \new_Sorter100|15753_  = \new_Sorter100|15653_  & \new_Sorter100|15654_ ;
  assign \new_Sorter100|15754_  = \new_Sorter100|15653_  | \new_Sorter100|15654_ ;
  assign \new_Sorter100|15755_  = \new_Sorter100|15655_  & \new_Sorter100|15656_ ;
  assign \new_Sorter100|15756_  = \new_Sorter100|15655_  | \new_Sorter100|15656_ ;
  assign \new_Sorter100|15757_  = \new_Sorter100|15657_  & \new_Sorter100|15658_ ;
  assign \new_Sorter100|15758_  = \new_Sorter100|15657_  | \new_Sorter100|15658_ ;
  assign \new_Sorter100|15759_  = \new_Sorter100|15659_  & \new_Sorter100|15660_ ;
  assign \new_Sorter100|15760_  = \new_Sorter100|15659_  | \new_Sorter100|15660_ ;
  assign \new_Sorter100|15761_  = \new_Sorter100|15661_  & \new_Sorter100|15662_ ;
  assign \new_Sorter100|15762_  = \new_Sorter100|15661_  | \new_Sorter100|15662_ ;
  assign \new_Sorter100|15763_  = \new_Sorter100|15663_  & \new_Sorter100|15664_ ;
  assign \new_Sorter100|15764_  = \new_Sorter100|15663_  | \new_Sorter100|15664_ ;
  assign \new_Sorter100|15765_  = \new_Sorter100|15665_  & \new_Sorter100|15666_ ;
  assign \new_Sorter100|15766_  = \new_Sorter100|15665_  | \new_Sorter100|15666_ ;
  assign \new_Sorter100|15767_  = \new_Sorter100|15667_  & \new_Sorter100|15668_ ;
  assign \new_Sorter100|15768_  = \new_Sorter100|15667_  | \new_Sorter100|15668_ ;
  assign \new_Sorter100|15769_  = \new_Sorter100|15669_  & \new_Sorter100|15670_ ;
  assign \new_Sorter100|15770_  = \new_Sorter100|15669_  | \new_Sorter100|15670_ ;
  assign \new_Sorter100|15771_  = \new_Sorter100|15671_  & \new_Sorter100|15672_ ;
  assign \new_Sorter100|15772_  = \new_Sorter100|15671_  | \new_Sorter100|15672_ ;
  assign \new_Sorter100|15773_  = \new_Sorter100|15673_  & \new_Sorter100|15674_ ;
  assign \new_Sorter100|15774_  = \new_Sorter100|15673_  | \new_Sorter100|15674_ ;
  assign \new_Sorter100|15775_  = \new_Sorter100|15675_  & \new_Sorter100|15676_ ;
  assign \new_Sorter100|15776_  = \new_Sorter100|15675_  | \new_Sorter100|15676_ ;
  assign \new_Sorter100|15777_  = \new_Sorter100|15677_  & \new_Sorter100|15678_ ;
  assign \new_Sorter100|15778_  = \new_Sorter100|15677_  | \new_Sorter100|15678_ ;
  assign \new_Sorter100|15779_  = \new_Sorter100|15679_  & \new_Sorter100|15680_ ;
  assign \new_Sorter100|15780_  = \new_Sorter100|15679_  | \new_Sorter100|15680_ ;
  assign \new_Sorter100|15781_  = \new_Sorter100|15681_  & \new_Sorter100|15682_ ;
  assign \new_Sorter100|15782_  = \new_Sorter100|15681_  | \new_Sorter100|15682_ ;
  assign \new_Sorter100|15783_  = \new_Sorter100|15683_  & \new_Sorter100|15684_ ;
  assign \new_Sorter100|15784_  = \new_Sorter100|15683_  | \new_Sorter100|15684_ ;
  assign \new_Sorter100|15785_  = \new_Sorter100|15685_  & \new_Sorter100|15686_ ;
  assign \new_Sorter100|15786_  = \new_Sorter100|15685_  | \new_Sorter100|15686_ ;
  assign \new_Sorter100|15787_  = \new_Sorter100|15687_  & \new_Sorter100|15688_ ;
  assign \new_Sorter100|15788_  = \new_Sorter100|15687_  | \new_Sorter100|15688_ ;
  assign \new_Sorter100|15789_  = \new_Sorter100|15689_  & \new_Sorter100|15690_ ;
  assign \new_Sorter100|15790_  = \new_Sorter100|15689_  | \new_Sorter100|15690_ ;
  assign \new_Sorter100|15791_  = \new_Sorter100|15691_  & \new_Sorter100|15692_ ;
  assign \new_Sorter100|15792_  = \new_Sorter100|15691_  | \new_Sorter100|15692_ ;
  assign \new_Sorter100|15793_  = \new_Sorter100|15693_  & \new_Sorter100|15694_ ;
  assign \new_Sorter100|15794_  = \new_Sorter100|15693_  | \new_Sorter100|15694_ ;
  assign \new_Sorter100|15795_  = \new_Sorter100|15695_  & \new_Sorter100|15696_ ;
  assign \new_Sorter100|15796_  = \new_Sorter100|15695_  | \new_Sorter100|15696_ ;
  assign \new_Sorter100|15797_  = \new_Sorter100|15697_  & \new_Sorter100|15698_ ;
  assign \new_Sorter100|15798_  = \new_Sorter100|15697_  | \new_Sorter100|15698_ ;
  assign \new_Sorter100|15800_  = \new_Sorter100|15700_  & \new_Sorter100|15701_ ;
  assign \new_Sorter100|15801_  = \new_Sorter100|15700_  | \new_Sorter100|15701_ ;
  assign \new_Sorter100|15802_  = \new_Sorter100|15702_  & \new_Sorter100|15703_ ;
  assign \new_Sorter100|15803_  = \new_Sorter100|15702_  | \new_Sorter100|15703_ ;
  assign \new_Sorter100|15804_  = \new_Sorter100|15704_  & \new_Sorter100|15705_ ;
  assign \new_Sorter100|15805_  = \new_Sorter100|15704_  | \new_Sorter100|15705_ ;
  assign \new_Sorter100|15806_  = \new_Sorter100|15706_  & \new_Sorter100|15707_ ;
  assign \new_Sorter100|15807_  = \new_Sorter100|15706_  | \new_Sorter100|15707_ ;
  assign \new_Sorter100|15808_  = \new_Sorter100|15708_  & \new_Sorter100|15709_ ;
  assign \new_Sorter100|15809_  = \new_Sorter100|15708_  | \new_Sorter100|15709_ ;
  assign \new_Sorter100|15810_  = \new_Sorter100|15710_  & \new_Sorter100|15711_ ;
  assign \new_Sorter100|15811_  = \new_Sorter100|15710_  | \new_Sorter100|15711_ ;
  assign \new_Sorter100|15812_  = \new_Sorter100|15712_  & \new_Sorter100|15713_ ;
  assign \new_Sorter100|15813_  = \new_Sorter100|15712_  | \new_Sorter100|15713_ ;
  assign \new_Sorter100|15814_  = \new_Sorter100|15714_  & \new_Sorter100|15715_ ;
  assign \new_Sorter100|15815_  = \new_Sorter100|15714_  | \new_Sorter100|15715_ ;
  assign \new_Sorter100|15816_  = \new_Sorter100|15716_  & \new_Sorter100|15717_ ;
  assign \new_Sorter100|15817_  = \new_Sorter100|15716_  | \new_Sorter100|15717_ ;
  assign \new_Sorter100|15818_  = \new_Sorter100|15718_  & \new_Sorter100|15719_ ;
  assign \new_Sorter100|15819_  = \new_Sorter100|15718_  | \new_Sorter100|15719_ ;
  assign \new_Sorter100|15820_  = \new_Sorter100|15720_  & \new_Sorter100|15721_ ;
  assign \new_Sorter100|15821_  = \new_Sorter100|15720_  | \new_Sorter100|15721_ ;
  assign \new_Sorter100|15822_  = \new_Sorter100|15722_  & \new_Sorter100|15723_ ;
  assign \new_Sorter100|15823_  = \new_Sorter100|15722_  | \new_Sorter100|15723_ ;
  assign \new_Sorter100|15824_  = \new_Sorter100|15724_  & \new_Sorter100|15725_ ;
  assign \new_Sorter100|15825_  = \new_Sorter100|15724_  | \new_Sorter100|15725_ ;
  assign \new_Sorter100|15826_  = \new_Sorter100|15726_  & \new_Sorter100|15727_ ;
  assign \new_Sorter100|15827_  = \new_Sorter100|15726_  | \new_Sorter100|15727_ ;
  assign \new_Sorter100|15828_  = \new_Sorter100|15728_  & \new_Sorter100|15729_ ;
  assign \new_Sorter100|15829_  = \new_Sorter100|15728_  | \new_Sorter100|15729_ ;
  assign \new_Sorter100|15830_  = \new_Sorter100|15730_  & \new_Sorter100|15731_ ;
  assign \new_Sorter100|15831_  = \new_Sorter100|15730_  | \new_Sorter100|15731_ ;
  assign \new_Sorter100|15832_  = \new_Sorter100|15732_  & \new_Sorter100|15733_ ;
  assign \new_Sorter100|15833_  = \new_Sorter100|15732_  | \new_Sorter100|15733_ ;
  assign \new_Sorter100|15834_  = \new_Sorter100|15734_  & \new_Sorter100|15735_ ;
  assign \new_Sorter100|15835_  = \new_Sorter100|15734_  | \new_Sorter100|15735_ ;
  assign \new_Sorter100|15836_  = \new_Sorter100|15736_  & \new_Sorter100|15737_ ;
  assign \new_Sorter100|15837_  = \new_Sorter100|15736_  | \new_Sorter100|15737_ ;
  assign \new_Sorter100|15838_  = \new_Sorter100|15738_  & \new_Sorter100|15739_ ;
  assign \new_Sorter100|15839_  = \new_Sorter100|15738_  | \new_Sorter100|15739_ ;
  assign \new_Sorter100|15840_  = \new_Sorter100|15740_  & \new_Sorter100|15741_ ;
  assign \new_Sorter100|15841_  = \new_Sorter100|15740_  | \new_Sorter100|15741_ ;
  assign \new_Sorter100|15842_  = \new_Sorter100|15742_  & \new_Sorter100|15743_ ;
  assign \new_Sorter100|15843_  = \new_Sorter100|15742_  | \new_Sorter100|15743_ ;
  assign \new_Sorter100|15844_  = \new_Sorter100|15744_  & \new_Sorter100|15745_ ;
  assign \new_Sorter100|15845_  = \new_Sorter100|15744_  | \new_Sorter100|15745_ ;
  assign \new_Sorter100|15846_  = \new_Sorter100|15746_  & \new_Sorter100|15747_ ;
  assign \new_Sorter100|15847_  = \new_Sorter100|15746_  | \new_Sorter100|15747_ ;
  assign \new_Sorter100|15848_  = \new_Sorter100|15748_  & \new_Sorter100|15749_ ;
  assign \new_Sorter100|15849_  = \new_Sorter100|15748_  | \new_Sorter100|15749_ ;
  assign \new_Sorter100|15850_  = \new_Sorter100|15750_  & \new_Sorter100|15751_ ;
  assign \new_Sorter100|15851_  = \new_Sorter100|15750_  | \new_Sorter100|15751_ ;
  assign \new_Sorter100|15852_  = \new_Sorter100|15752_  & \new_Sorter100|15753_ ;
  assign \new_Sorter100|15853_  = \new_Sorter100|15752_  | \new_Sorter100|15753_ ;
  assign \new_Sorter100|15854_  = \new_Sorter100|15754_  & \new_Sorter100|15755_ ;
  assign \new_Sorter100|15855_  = \new_Sorter100|15754_  | \new_Sorter100|15755_ ;
  assign \new_Sorter100|15856_  = \new_Sorter100|15756_  & \new_Sorter100|15757_ ;
  assign \new_Sorter100|15857_  = \new_Sorter100|15756_  | \new_Sorter100|15757_ ;
  assign \new_Sorter100|15858_  = \new_Sorter100|15758_  & \new_Sorter100|15759_ ;
  assign \new_Sorter100|15859_  = \new_Sorter100|15758_  | \new_Sorter100|15759_ ;
  assign \new_Sorter100|15860_  = \new_Sorter100|15760_  & \new_Sorter100|15761_ ;
  assign \new_Sorter100|15861_  = \new_Sorter100|15760_  | \new_Sorter100|15761_ ;
  assign \new_Sorter100|15862_  = \new_Sorter100|15762_  & \new_Sorter100|15763_ ;
  assign \new_Sorter100|15863_  = \new_Sorter100|15762_  | \new_Sorter100|15763_ ;
  assign \new_Sorter100|15864_  = \new_Sorter100|15764_  & \new_Sorter100|15765_ ;
  assign \new_Sorter100|15865_  = \new_Sorter100|15764_  | \new_Sorter100|15765_ ;
  assign \new_Sorter100|15866_  = \new_Sorter100|15766_  & \new_Sorter100|15767_ ;
  assign \new_Sorter100|15867_  = \new_Sorter100|15766_  | \new_Sorter100|15767_ ;
  assign \new_Sorter100|15868_  = \new_Sorter100|15768_  & \new_Sorter100|15769_ ;
  assign \new_Sorter100|15869_  = \new_Sorter100|15768_  | \new_Sorter100|15769_ ;
  assign \new_Sorter100|15870_  = \new_Sorter100|15770_  & \new_Sorter100|15771_ ;
  assign \new_Sorter100|15871_  = \new_Sorter100|15770_  | \new_Sorter100|15771_ ;
  assign \new_Sorter100|15872_  = \new_Sorter100|15772_  & \new_Sorter100|15773_ ;
  assign \new_Sorter100|15873_  = \new_Sorter100|15772_  | \new_Sorter100|15773_ ;
  assign \new_Sorter100|15874_  = \new_Sorter100|15774_  & \new_Sorter100|15775_ ;
  assign \new_Sorter100|15875_  = \new_Sorter100|15774_  | \new_Sorter100|15775_ ;
  assign \new_Sorter100|15876_  = \new_Sorter100|15776_  & \new_Sorter100|15777_ ;
  assign \new_Sorter100|15877_  = \new_Sorter100|15776_  | \new_Sorter100|15777_ ;
  assign \new_Sorter100|15878_  = \new_Sorter100|15778_  & \new_Sorter100|15779_ ;
  assign \new_Sorter100|15879_  = \new_Sorter100|15778_  | \new_Sorter100|15779_ ;
  assign \new_Sorter100|15880_  = \new_Sorter100|15780_  & \new_Sorter100|15781_ ;
  assign \new_Sorter100|15881_  = \new_Sorter100|15780_  | \new_Sorter100|15781_ ;
  assign \new_Sorter100|15882_  = \new_Sorter100|15782_  & \new_Sorter100|15783_ ;
  assign \new_Sorter100|15883_  = \new_Sorter100|15782_  | \new_Sorter100|15783_ ;
  assign \new_Sorter100|15884_  = \new_Sorter100|15784_  & \new_Sorter100|15785_ ;
  assign \new_Sorter100|15885_  = \new_Sorter100|15784_  | \new_Sorter100|15785_ ;
  assign \new_Sorter100|15886_  = \new_Sorter100|15786_  & \new_Sorter100|15787_ ;
  assign \new_Sorter100|15887_  = \new_Sorter100|15786_  | \new_Sorter100|15787_ ;
  assign \new_Sorter100|15888_  = \new_Sorter100|15788_  & \new_Sorter100|15789_ ;
  assign \new_Sorter100|15889_  = \new_Sorter100|15788_  | \new_Sorter100|15789_ ;
  assign \new_Sorter100|15890_  = \new_Sorter100|15790_  & \new_Sorter100|15791_ ;
  assign \new_Sorter100|15891_  = \new_Sorter100|15790_  | \new_Sorter100|15791_ ;
  assign \new_Sorter100|15892_  = \new_Sorter100|15792_  & \new_Sorter100|15793_ ;
  assign \new_Sorter100|15893_  = \new_Sorter100|15792_  | \new_Sorter100|15793_ ;
  assign \new_Sorter100|15894_  = \new_Sorter100|15794_  & \new_Sorter100|15795_ ;
  assign \new_Sorter100|15895_  = \new_Sorter100|15794_  | \new_Sorter100|15795_ ;
  assign \new_Sorter100|15896_  = \new_Sorter100|15796_  & \new_Sorter100|15797_ ;
  assign \new_Sorter100|15897_  = \new_Sorter100|15796_  | \new_Sorter100|15797_ ;
  assign \new_Sorter100|15898_  = \new_Sorter100|15798_  & \new_Sorter100|15799_ ;
  assign \new_Sorter100|15899_  = \new_Sorter100|15798_  | \new_Sorter100|15799_ ;
  assign \new_Sorter100|15900_  = \new_Sorter100|15800_ ;
  assign \new_Sorter100|15999_  = \new_Sorter100|15899_ ;
  assign \new_Sorter100|15901_  = \new_Sorter100|15801_  & \new_Sorter100|15802_ ;
  assign \new_Sorter100|15902_  = \new_Sorter100|15801_  | \new_Sorter100|15802_ ;
  assign \new_Sorter100|15903_  = \new_Sorter100|15803_  & \new_Sorter100|15804_ ;
  assign \new_Sorter100|15904_  = \new_Sorter100|15803_  | \new_Sorter100|15804_ ;
  assign \new_Sorter100|15905_  = \new_Sorter100|15805_  & \new_Sorter100|15806_ ;
  assign \new_Sorter100|15906_  = \new_Sorter100|15805_  | \new_Sorter100|15806_ ;
  assign \new_Sorter100|15907_  = \new_Sorter100|15807_  & \new_Sorter100|15808_ ;
  assign \new_Sorter100|15908_  = \new_Sorter100|15807_  | \new_Sorter100|15808_ ;
  assign \new_Sorter100|15909_  = \new_Sorter100|15809_  & \new_Sorter100|15810_ ;
  assign \new_Sorter100|15910_  = \new_Sorter100|15809_  | \new_Sorter100|15810_ ;
  assign \new_Sorter100|15911_  = \new_Sorter100|15811_  & \new_Sorter100|15812_ ;
  assign \new_Sorter100|15912_  = \new_Sorter100|15811_  | \new_Sorter100|15812_ ;
  assign \new_Sorter100|15913_  = \new_Sorter100|15813_  & \new_Sorter100|15814_ ;
  assign \new_Sorter100|15914_  = \new_Sorter100|15813_  | \new_Sorter100|15814_ ;
  assign \new_Sorter100|15915_  = \new_Sorter100|15815_  & \new_Sorter100|15816_ ;
  assign \new_Sorter100|15916_  = \new_Sorter100|15815_  | \new_Sorter100|15816_ ;
  assign \new_Sorter100|15917_  = \new_Sorter100|15817_  & \new_Sorter100|15818_ ;
  assign \new_Sorter100|15918_  = \new_Sorter100|15817_  | \new_Sorter100|15818_ ;
  assign \new_Sorter100|15919_  = \new_Sorter100|15819_  & \new_Sorter100|15820_ ;
  assign \new_Sorter100|15920_  = \new_Sorter100|15819_  | \new_Sorter100|15820_ ;
  assign \new_Sorter100|15921_  = \new_Sorter100|15821_  & \new_Sorter100|15822_ ;
  assign \new_Sorter100|15922_  = \new_Sorter100|15821_  | \new_Sorter100|15822_ ;
  assign \new_Sorter100|15923_  = \new_Sorter100|15823_  & \new_Sorter100|15824_ ;
  assign \new_Sorter100|15924_  = \new_Sorter100|15823_  | \new_Sorter100|15824_ ;
  assign \new_Sorter100|15925_  = \new_Sorter100|15825_  & \new_Sorter100|15826_ ;
  assign \new_Sorter100|15926_  = \new_Sorter100|15825_  | \new_Sorter100|15826_ ;
  assign \new_Sorter100|15927_  = \new_Sorter100|15827_  & \new_Sorter100|15828_ ;
  assign \new_Sorter100|15928_  = \new_Sorter100|15827_  | \new_Sorter100|15828_ ;
  assign \new_Sorter100|15929_  = \new_Sorter100|15829_  & \new_Sorter100|15830_ ;
  assign \new_Sorter100|15930_  = \new_Sorter100|15829_  | \new_Sorter100|15830_ ;
  assign \new_Sorter100|15931_  = \new_Sorter100|15831_  & \new_Sorter100|15832_ ;
  assign \new_Sorter100|15932_  = \new_Sorter100|15831_  | \new_Sorter100|15832_ ;
  assign \new_Sorter100|15933_  = \new_Sorter100|15833_  & \new_Sorter100|15834_ ;
  assign \new_Sorter100|15934_  = \new_Sorter100|15833_  | \new_Sorter100|15834_ ;
  assign \new_Sorter100|15935_  = \new_Sorter100|15835_  & \new_Sorter100|15836_ ;
  assign \new_Sorter100|15936_  = \new_Sorter100|15835_  | \new_Sorter100|15836_ ;
  assign \new_Sorter100|15937_  = \new_Sorter100|15837_  & \new_Sorter100|15838_ ;
  assign \new_Sorter100|15938_  = \new_Sorter100|15837_  | \new_Sorter100|15838_ ;
  assign \new_Sorter100|15939_  = \new_Sorter100|15839_  & \new_Sorter100|15840_ ;
  assign \new_Sorter100|15940_  = \new_Sorter100|15839_  | \new_Sorter100|15840_ ;
  assign \new_Sorter100|15941_  = \new_Sorter100|15841_  & \new_Sorter100|15842_ ;
  assign \new_Sorter100|15942_  = \new_Sorter100|15841_  | \new_Sorter100|15842_ ;
  assign \new_Sorter100|15943_  = \new_Sorter100|15843_  & \new_Sorter100|15844_ ;
  assign \new_Sorter100|15944_  = \new_Sorter100|15843_  | \new_Sorter100|15844_ ;
  assign \new_Sorter100|15945_  = \new_Sorter100|15845_  & \new_Sorter100|15846_ ;
  assign \new_Sorter100|15946_  = \new_Sorter100|15845_  | \new_Sorter100|15846_ ;
  assign \new_Sorter100|15947_  = \new_Sorter100|15847_  & \new_Sorter100|15848_ ;
  assign \new_Sorter100|15948_  = \new_Sorter100|15847_  | \new_Sorter100|15848_ ;
  assign \new_Sorter100|15949_  = \new_Sorter100|15849_  & \new_Sorter100|15850_ ;
  assign \new_Sorter100|15950_  = \new_Sorter100|15849_  | \new_Sorter100|15850_ ;
  assign \new_Sorter100|15951_  = \new_Sorter100|15851_  & \new_Sorter100|15852_ ;
  assign \new_Sorter100|15952_  = \new_Sorter100|15851_  | \new_Sorter100|15852_ ;
  assign \new_Sorter100|15953_  = \new_Sorter100|15853_  & \new_Sorter100|15854_ ;
  assign \new_Sorter100|15954_  = \new_Sorter100|15853_  | \new_Sorter100|15854_ ;
  assign \new_Sorter100|15955_  = \new_Sorter100|15855_  & \new_Sorter100|15856_ ;
  assign \new_Sorter100|15956_  = \new_Sorter100|15855_  | \new_Sorter100|15856_ ;
  assign \new_Sorter100|15957_  = \new_Sorter100|15857_  & \new_Sorter100|15858_ ;
  assign \new_Sorter100|15958_  = \new_Sorter100|15857_  | \new_Sorter100|15858_ ;
  assign \new_Sorter100|15959_  = \new_Sorter100|15859_  & \new_Sorter100|15860_ ;
  assign \new_Sorter100|15960_  = \new_Sorter100|15859_  | \new_Sorter100|15860_ ;
  assign \new_Sorter100|15961_  = \new_Sorter100|15861_  & \new_Sorter100|15862_ ;
  assign \new_Sorter100|15962_  = \new_Sorter100|15861_  | \new_Sorter100|15862_ ;
  assign \new_Sorter100|15963_  = \new_Sorter100|15863_  & \new_Sorter100|15864_ ;
  assign \new_Sorter100|15964_  = \new_Sorter100|15863_  | \new_Sorter100|15864_ ;
  assign \new_Sorter100|15965_  = \new_Sorter100|15865_  & \new_Sorter100|15866_ ;
  assign \new_Sorter100|15966_  = \new_Sorter100|15865_  | \new_Sorter100|15866_ ;
  assign \new_Sorter100|15967_  = \new_Sorter100|15867_  & \new_Sorter100|15868_ ;
  assign \new_Sorter100|15968_  = \new_Sorter100|15867_  | \new_Sorter100|15868_ ;
  assign \new_Sorter100|15969_  = \new_Sorter100|15869_  & \new_Sorter100|15870_ ;
  assign \new_Sorter100|15970_  = \new_Sorter100|15869_  | \new_Sorter100|15870_ ;
  assign \new_Sorter100|15971_  = \new_Sorter100|15871_  & \new_Sorter100|15872_ ;
  assign \new_Sorter100|15972_  = \new_Sorter100|15871_  | \new_Sorter100|15872_ ;
  assign \new_Sorter100|15973_  = \new_Sorter100|15873_  & \new_Sorter100|15874_ ;
  assign \new_Sorter100|15974_  = \new_Sorter100|15873_  | \new_Sorter100|15874_ ;
  assign \new_Sorter100|15975_  = \new_Sorter100|15875_  & \new_Sorter100|15876_ ;
  assign \new_Sorter100|15976_  = \new_Sorter100|15875_  | \new_Sorter100|15876_ ;
  assign \new_Sorter100|15977_  = \new_Sorter100|15877_  & \new_Sorter100|15878_ ;
  assign \new_Sorter100|15978_  = \new_Sorter100|15877_  | \new_Sorter100|15878_ ;
  assign \new_Sorter100|15979_  = \new_Sorter100|15879_  & \new_Sorter100|15880_ ;
  assign \new_Sorter100|15980_  = \new_Sorter100|15879_  | \new_Sorter100|15880_ ;
  assign \new_Sorter100|15981_  = \new_Sorter100|15881_  & \new_Sorter100|15882_ ;
  assign \new_Sorter100|15982_  = \new_Sorter100|15881_  | \new_Sorter100|15882_ ;
  assign \new_Sorter100|15983_  = \new_Sorter100|15883_  & \new_Sorter100|15884_ ;
  assign \new_Sorter100|15984_  = \new_Sorter100|15883_  | \new_Sorter100|15884_ ;
  assign \new_Sorter100|15985_  = \new_Sorter100|15885_  & \new_Sorter100|15886_ ;
  assign \new_Sorter100|15986_  = \new_Sorter100|15885_  | \new_Sorter100|15886_ ;
  assign \new_Sorter100|15987_  = \new_Sorter100|15887_  & \new_Sorter100|15888_ ;
  assign \new_Sorter100|15988_  = \new_Sorter100|15887_  | \new_Sorter100|15888_ ;
  assign \new_Sorter100|15989_  = \new_Sorter100|15889_  & \new_Sorter100|15890_ ;
  assign \new_Sorter100|15990_  = \new_Sorter100|15889_  | \new_Sorter100|15890_ ;
  assign \new_Sorter100|15991_  = \new_Sorter100|15891_  & \new_Sorter100|15892_ ;
  assign \new_Sorter100|15992_  = \new_Sorter100|15891_  | \new_Sorter100|15892_ ;
  assign \new_Sorter100|15993_  = \new_Sorter100|15893_  & \new_Sorter100|15894_ ;
  assign \new_Sorter100|15994_  = \new_Sorter100|15893_  | \new_Sorter100|15894_ ;
  assign \new_Sorter100|15995_  = \new_Sorter100|15895_  & \new_Sorter100|15896_ ;
  assign \new_Sorter100|15996_  = \new_Sorter100|15895_  | \new_Sorter100|15896_ ;
  assign \new_Sorter100|15997_  = \new_Sorter100|15897_  & \new_Sorter100|15898_ ;
  assign \new_Sorter100|15998_  = \new_Sorter100|15897_  | \new_Sorter100|15898_ ;
  assign \new_Sorter100|16000_  = \new_Sorter100|15900_  & \new_Sorter100|15901_ ;
  assign \new_Sorter100|16001_  = \new_Sorter100|15900_  | \new_Sorter100|15901_ ;
  assign \new_Sorter100|16002_  = \new_Sorter100|15902_  & \new_Sorter100|15903_ ;
  assign \new_Sorter100|16003_  = \new_Sorter100|15902_  | \new_Sorter100|15903_ ;
  assign \new_Sorter100|16004_  = \new_Sorter100|15904_  & \new_Sorter100|15905_ ;
  assign \new_Sorter100|16005_  = \new_Sorter100|15904_  | \new_Sorter100|15905_ ;
  assign \new_Sorter100|16006_  = \new_Sorter100|15906_  & \new_Sorter100|15907_ ;
  assign \new_Sorter100|16007_  = \new_Sorter100|15906_  | \new_Sorter100|15907_ ;
  assign \new_Sorter100|16008_  = \new_Sorter100|15908_  & \new_Sorter100|15909_ ;
  assign \new_Sorter100|16009_  = \new_Sorter100|15908_  | \new_Sorter100|15909_ ;
  assign \new_Sorter100|16010_  = \new_Sorter100|15910_  & \new_Sorter100|15911_ ;
  assign \new_Sorter100|16011_  = \new_Sorter100|15910_  | \new_Sorter100|15911_ ;
  assign \new_Sorter100|16012_  = \new_Sorter100|15912_  & \new_Sorter100|15913_ ;
  assign \new_Sorter100|16013_  = \new_Sorter100|15912_  | \new_Sorter100|15913_ ;
  assign \new_Sorter100|16014_  = \new_Sorter100|15914_  & \new_Sorter100|15915_ ;
  assign \new_Sorter100|16015_  = \new_Sorter100|15914_  | \new_Sorter100|15915_ ;
  assign \new_Sorter100|16016_  = \new_Sorter100|15916_  & \new_Sorter100|15917_ ;
  assign \new_Sorter100|16017_  = \new_Sorter100|15916_  | \new_Sorter100|15917_ ;
  assign \new_Sorter100|16018_  = \new_Sorter100|15918_  & \new_Sorter100|15919_ ;
  assign \new_Sorter100|16019_  = \new_Sorter100|15918_  | \new_Sorter100|15919_ ;
  assign \new_Sorter100|16020_  = \new_Sorter100|15920_  & \new_Sorter100|15921_ ;
  assign \new_Sorter100|16021_  = \new_Sorter100|15920_  | \new_Sorter100|15921_ ;
  assign \new_Sorter100|16022_  = \new_Sorter100|15922_  & \new_Sorter100|15923_ ;
  assign \new_Sorter100|16023_  = \new_Sorter100|15922_  | \new_Sorter100|15923_ ;
  assign \new_Sorter100|16024_  = \new_Sorter100|15924_  & \new_Sorter100|15925_ ;
  assign \new_Sorter100|16025_  = \new_Sorter100|15924_  | \new_Sorter100|15925_ ;
  assign \new_Sorter100|16026_  = \new_Sorter100|15926_  & \new_Sorter100|15927_ ;
  assign \new_Sorter100|16027_  = \new_Sorter100|15926_  | \new_Sorter100|15927_ ;
  assign \new_Sorter100|16028_  = \new_Sorter100|15928_  & \new_Sorter100|15929_ ;
  assign \new_Sorter100|16029_  = \new_Sorter100|15928_  | \new_Sorter100|15929_ ;
  assign \new_Sorter100|16030_  = \new_Sorter100|15930_  & \new_Sorter100|15931_ ;
  assign \new_Sorter100|16031_  = \new_Sorter100|15930_  | \new_Sorter100|15931_ ;
  assign \new_Sorter100|16032_  = \new_Sorter100|15932_  & \new_Sorter100|15933_ ;
  assign \new_Sorter100|16033_  = \new_Sorter100|15932_  | \new_Sorter100|15933_ ;
  assign \new_Sorter100|16034_  = \new_Sorter100|15934_  & \new_Sorter100|15935_ ;
  assign \new_Sorter100|16035_  = \new_Sorter100|15934_  | \new_Sorter100|15935_ ;
  assign \new_Sorter100|16036_  = \new_Sorter100|15936_  & \new_Sorter100|15937_ ;
  assign \new_Sorter100|16037_  = \new_Sorter100|15936_  | \new_Sorter100|15937_ ;
  assign \new_Sorter100|16038_  = \new_Sorter100|15938_  & \new_Sorter100|15939_ ;
  assign \new_Sorter100|16039_  = \new_Sorter100|15938_  | \new_Sorter100|15939_ ;
  assign \new_Sorter100|16040_  = \new_Sorter100|15940_  & \new_Sorter100|15941_ ;
  assign \new_Sorter100|16041_  = \new_Sorter100|15940_  | \new_Sorter100|15941_ ;
  assign \new_Sorter100|16042_  = \new_Sorter100|15942_  & \new_Sorter100|15943_ ;
  assign \new_Sorter100|16043_  = \new_Sorter100|15942_  | \new_Sorter100|15943_ ;
  assign \new_Sorter100|16044_  = \new_Sorter100|15944_  & \new_Sorter100|15945_ ;
  assign \new_Sorter100|16045_  = \new_Sorter100|15944_  | \new_Sorter100|15945_ ;
  assign \new_Sorter100|16046_  = \new_Sorter100|15946_  & \new_Sorter100|15947_ ;
  assign \new_Sorter100|16047_  = \new_Sorter100|15946_  | \new_Sorter100|15947_ ;
  assign \new_Sorter100|16048_  = \new_Sorter100|15948_  & \new_Sorter100|15949_ ;
  assign \new_Sorter100|16049_  = \new_Sorter100|15948_  | \new_Sorter100|15949_ ;
  assign \new_Sorter100|16050_  = \new_Sorter100|15950_  & \new_Sorter100|15951_ ;
  assign \new_Sorter100|16051_  = \new_Sorter100|15950_  | \new_Sorter100|15951_ ;
  assign \new_Sorter100|16052_  = \new_Sorter100|15952_  & \new_Sorter100|15953_ ;
  assign \new_Sorter100|16053_  = \new_Sorter100|15952_  | \new_Sorter100|15953_ ;
  assign \new_Sorter100|16054_  = \new_Sorter100|15954_  & \new_Sorter100|15955_ ;
  assign \new_Sorter100|16055_  = \new_Sorter100|15954_  | \new_Sorter100|15955_ ;
  assign \new_Sorter100|16056_  = \new_Sorter100|15956_  & \new_Sorter100|15957_ ;
  assign \new_Sorter100|16057_  = \new_Sorter100|15956_  | \new_Sorter100|15957_ ;
  assign \new_Sorter100|16058_  = \new_Sorter100|15958_  & \new_Sorter100|15959_ ;
  assign \new_Sorter100|16059_  = \new_Sorter100|15958_  | \new_Sorter100|15959_ ;
  assign \new_Sorter100|16060_  = \new_Sorter100|15960_  & \new_Sorter100|15961_ ;
  assign \new_Sorter100|16061_  = \new_Sorter100|15960_  | \new_Sorter100|15961_ ;
  assign \new_Sorter100|16062_  = \new_Sorter100|15962_  & \new_Sorter100|15963_ ;
  assign \new_Sorter100|16063_  = \new_Sorter100|15962_  | \new_Sorter100|15963_ ;
  assign \new_Sorter100|16064_  = \new_Sorter100|15964_  & \new_Sorter100|15965_ ;
  assign \new_Sorter100|16065_  = \new_Sorter100|15964_  | \new_Sorter100|15965_ ;
  assign \new_Sorter100|16066_  = \new_Sorter100|15966_  & \new_Sorter100|15967_ ;
  assign \new_Sorter100|16067_  = \new_Sorter100|15966_  | \new_Sorter100|15967_ ;
  assign \new_Sorter100|16068_  = \new_Sorter100|15968_  & \new_Sorter100|15969_ ;
  assign \new_Sorter100|16069_  = \new_Sorter100|15968_  | \new_Sorter100|15969_ ;
  assign \new_Sorter100|16070_  = \new_Sorter100|15970_  & \new_Sorter100|15971_ ;
  assign \new_Sorter100|16071_  = \new_Sorter100|15970_  | \new_Sorter100|15971_ ;
  assign \new_Sorter100|16072_  = \new_Sorter100|15972_  & \new_Sorter100|15973_ ;
  assign \new_Sorter100|16073_  = \new_Sorter100|15972_  | \new_Sorter100|15973_ ;
  assign \new_Sorter100|16074_  = \new_Sorter100|15974_  & \new_Sorter100|15975_ ;
  assign \new_Sorter100|16075_  = \new_Sorter100|15974_  | \new_Sorter100|15975_ ;
  assign \new_Sorter100|16076_  = \new_Sorter100|15976_  & \new_Sorter100|15977_ ;
  assign \new_Sorter100|16077_  = \new_Sorter100|15976_  | \new_Sorter100|15977_ ;
  assign \new_Sorter100|16078_  = \new_Sorter100|15978_  & \new_Sorter100|15979_ ;
  assign \new_Sorter100|16079_  = \new_Sorter100|15978_  | \new_Sorter100|15979_ ;
  assign \new_Sorter100|16080_  = \new_Sorter100|15980_  & \new_Sorter100|15981_ ;
  assign \new_Sorter100|16081_  = \new_Sorter100|15980_  | \new_Sorter100|15981_ ;
  assign \new_Sorter100|16082_  = \new_Sorter100|15982_  & \new_Sorter100|15983_ ;
  assign \new_Sorter100|16083_  = \new_Sorter100|15982_  | \new_Sorter100|15983_ ;
  assign \new_Sorter100|16084_  = \new_Sorter100|15984_  & \new_Sorter100|15985_ ;
  assign \new_Sorter100|16085_  = \new_Sorter100|15984_  | \new_Sorter100|15985_ ;
  assign \new_Sorter100|16086_  = \new_Sorter100|15986_  & \new_Sorter100|15987_ ;
  assign \new_Sorter100|16087_  = \new_Sorter100|15986_  | \new_Sorter100|15987_ ;
  assign \new_Sorter100|16088_  = \new_Sorter100|15988_  & \new_Sorter100|15989_ ;
  assign \new_Sorter100|16089_  = \new_Sorter100|15988_  | \new_Sorter100|15989_ ;
  assign \new_Sorter100|16090_  = \new_Sorter100|15990_  & \new_Sorter100|15991_ ;
  assign \new_Sorter100|16091_  = \new_Sorter100|15990_  | \new_Sorter100|15991_ ;
  assign \new_Sorter100|16092_  = \new_Sorter100|15992_  & \new_Sorter100|15993_ ;
  assign \new_Sorter100|16093_  = \new_Sorter100|15992_  | \new_Sorter100|15993_ ;
  assign \new_Sorter100|16094_  = \new_Sorter100|15994_  & \new_Sorter100|15995_ ;
  assign \new_Sorter100|16095_  = \new_Sorter100|15994_  | \new_Sorter100|15995_ ;
  assign \new_Sorter100|16096_  = \new_Sorter100|15996_  & \new_Sorter100|15997_ ;
  assign \new_Sorter100|16097_  = \new_Sorter100|15996_  | \new_Sorter100|15997_ ;
  assign \new_Sorter100|16098_  = \new_Sorter100|15998_  & \new_Sorter100|15999_ ;
  assign \new_Sorter100|16099_  = \new_Sorter100|15998_  | \new_Sorter100|15999_ ;
  assign \new_Sorter100|16100_  = \new_Sorter100|16000_ ;
  assign \new_Sorter100|16199_  = \new_Sorter100|16099_ ;
  assign \new_Sorter100|16101_  = \new_Sorter100|16001_  & \new_Sorter100|16002_ ;
  assign \new_Sorter100|16102_  = \new_Sorter100|16001_  | \new_Sorter100|16002_ ;
  assign \new_Sorter100|16103_  = \new_Sorter100|16003_  & \new_Sorter100|16004_ ;
  assign \new_Sorter100|16104_  = \new_Sorter100|16003_  | \new_Sorter100|16004_ ;
  assign \new_Sorter100|16105_  = \new_Sorter100|16005_  & \new_Sorter100|16006_ ;
  assign \new_Sorter100|16106_  = \new_Sorter100|16005_  | \new_Sorter100|16006_ ;
  assign \new_Sorter100|16107_  = \new_Sorter100|16007_  & \new_Sorter100|16008_ ;
  assign \new_Sorter100|16108_  = \new_Sorter100|16007_  | \new_Sorter100|16008_ ;
  assign \new_Sorter100|16109_  = \new_Sorter100|16009_  & \new_Sorter100|16010_ ;
  assign \new_Sorter100|16110_  = \new_Sorter100|16009_  | \new_Sorter100|16010_ ;
  assign \new_Sorter100|16111_  = \new_Sorter100|16011_  & \new_Sorter100|16012_ ;
  assign \new_Sorter100|16112_  = \new_Sorter100|16011_  | \new_Sorter100|16012_ ;
  assign \new_Sorter100|16113_  = \new_Sorter100|16013_  & \new_Sorter100|16014_ ;
  assign \new_Sorter100|16114_  = \new_Sorter100|16013_  | \new_Sorter100|16014_ ;
  assign \new_Sorter100|16115_  = \new_Sorter100|16015_  & \new_Sorter100|16016_ ;
  assign \new_Sorter100|16116_  = \new_Sorter100|16015_  | \new_Sorter100|16016_ ;
  assign \new_Sorter100|16117_  = \new_Sorter100|16017_  & \new_Sorter100|16018_ ;
  assign \new_Sorter100|16118_  = \new_Sorter100|16017_  | \new_Sorter100|16018_ ;
  assign \new_Sorter100|16119_  = \new_Sorter100|16019_  & \new_Sorter100|16020_ ;
  assign \new_Sorter100|16120_  = \new_Sorter100|16019_  | \new_Sorter100|16020_ ;
  assign \new_Sorter100|16121_  = \new_Sorter100|16021_  & \new_Sorter100|16022_ ;
  assign \new_Sorter100|16122_  = \new_Sorter100|16021_  | \new_Sorter100|16022_ ;
  assign \new_Sorter100|16123_  = \new_Sorter100|16023_  & \new_Sorter100|16024_ ;
  assign \new_Sorter100|16124_  = \new_Sorter100|16023_  | \new_Sorter100|16024_ ;
  assign \new_Sorter100|16125_  = \new_Sorter100|16025_  & \new_Sorter100|16026_ ;
  assign \new_Sorter100|16126_  = \new_Sorter100|16025_  | \new_Sorter100|16026_ ;
  assign \new_Sorter100|16127_  = \new_Sorter100|16027_  & \new_Sorter100|16028_ ;
  assign \new_Sorter100|16128_  = \new_Sorter100|16027_  | \new_Sorter100|16028_ ;
  assign \new_Sorter100|16129_  = \new_Sorter100|16029_  & \new_Sorter100|16030_ ;
  assign \new_Sorter100|16130_  = \new_Sorter100|16029_  | \new_Sorter100|16030_ ;
  assign \new_Sorter100|16131_  = \new_Sorter100|16031_  & \new_Sorter100|16032_ ;
  assign \new_Sorter100|16132_  = \new_Sorter100|16031_  | \new_Sorter100|16032_ ;
  assign \new_Sorter100|16133_  = \new_Sorter100|16033_  & \new_Sorter100|16034_ ;
  assign \new_Sorter100|16134_  = \new_Sorter100|16033_  | \new_Sorter100|16034_ ;
  assign \new_Sorter100|16135_  = \new_Sorter100|16035_  & \new_Sorter100|16036_ ;
  assign \new_Sorter100|16136_  = \new_Sorter100|16035_  | \new_Sorter100|16036_ ;
  assign \new_Sorter100|16137_  = \new_Sorter100|16037_  & \new_Sorter100|16038_ ;
  assign \new_Sorter100|16138_  = \new_Sorter100|16037_  | \new_Sorter100|16038_ ;
  assign \new_Sorter100|16139_  = \new_Sorter100|16039_  & \new_Sorter100|16040_ ;
  assign \new_Sorter100|16140_  = \new_Sorter100|16039_  | \new_Sorter100|16040_ ;
  assign \new_Sorter100|16141_  = \new_Sorter100|16041_  & \new_Sorter100|16042_ ;
  assign \new_Sorter100|16142_  = \new_Sorter100|16041_  | \new_Sorter100|16042_ ;
  assign \new_Sorter100|16143_  = \new_Sorter100|16043_  & \new_Sorter100|16044_ ;
  assign \new_Sorter100|16144_  = \new_Sorter100|16043_  | \new_Sorter100|16044_ ;
  assign \new_Sorter100|16145_  = \new_Sorter100|16045_  & \new_Sorter100|16046_ ;
  assign \new_Sorter100|16146_  = \new_Sorter100|16045_  | \new_Sorter100|16046_ ;
  assign \new_Sorter100|16147_  = \new_Sorter100|16047_  & \new_Sorter100|16048_ ;
  assign \new_Sorter100|16148_  = \new_Sorter100|16047_  | \new_Sorter100|16048_ ;
  assign \new_Sorter100|16149_  = \new_Sorter100|16049_  & \new_Sorter100|16050_ ;
  assign \new_Sorter100|16150_  = \new_Sorter100|16049_  | \new_Sorter100|16050_ ;
  assign \new_Sorter100|16151_  = \new_Sorter100|16051_  & \new_Sorter100|16052_ ;
  assign \new_Sorter100|16152_  = \new_Sorter100|16051_  | \new_Sorter100|16052_ ;
  assign \new_Sorter100|16153_  = \new_Sorter100|16053_  & \new_Sorter100|16054_ ;
  assign \new_Sorter100|16154_  = \new_Sorter100|16053_  | \new_Sorter100|16054_ ;
  assign \new_Sorter100|16155_  = \new_Sorter100|16055_  & \new_Sorter100|16056_ ;
  assign \new_Sorter100|16156_  = \new_Sorter100|16055_  | \new_Sorter100|16056_ ;
  assign \new_Sorter100|16157_  = \new_Sorter100|16057_  & \new_Sorter100|16058_ ;
  assign \new_Sorter100|16158_  = \new_Sorter100|16057_  | \new_Sorter100|16058_ ;
  assign \new_Sorter100|16159_  = \new_Sorter100|16059_  & \new_Sorter100|16060_ ;
  assign \new_Sorter100|16160_  = \new_Sorter100|16059_  | \new_Sorter100|16060_ ;
  assign \new_Sorter100|16161_  = \new_Sorter100|16061_  & \new_Sorter100|16062_ ;
  assign \new_Sorter100|16162_  = \new_Sorter100|16061_  | \new_Sorter100|16062_ ;
  assign \new_Sorter100|16163_  = \new_Sorter100|16063_  & \new_Sorter100|16064_ ;
  assign \new_Sorter100|16164_  = \new_Sorter100|16063_  | \new_Sorter100|16064_ ;
  assign \new_Sorter100|16165_  = \new_Sorter100|16065_  & \new_Sorter100|16066_ ;
  assign \new_Sorter100|16166_  = \new_Sorter100|16065_  | \new_Sorter100|16066_ ;
  assign \new_Sorter100|16167_  = \new_Sorter100|16067_  & \new_Sorter100|16068_ ;
  assign \new_Sorter100|16168_  = \new_Sorter100|16067_  | \new_Sorter100|16068_ ;
  assign \new_Sorter100|16169_  = \new_Sorter100|16069_  & \new_Sorter100|16070_ ;
  assign \new_Sorter100|16170_  = \new_Sorter100|16069_  | \new_Sorter100|16070_ ;
  assign \new_Sorter100|16171_  = \new_Sorter100|16071_  & \new_Sorter100|16072_ ;
  assign \new_Sorter100|16172_  = \new_Sorter100|16071_  | \new_Sorter100|16072_ ;
  assign \new_Sorter100|16173_  = \new_Sorter100|16073_  & \new_Sorter100|16074_ ;
  assign \new_Sorter100|16174_  = \new_Sorter100|16073_  | \new_Sorter100|16074_ ;
  assign \new_Sorter100|16175_  = \new_Sorter100|16075_  & \new_Sorter100|16076_ ;
  assign \new_Sorter100|16176_  = \new_Sorter100|16075_  | \new_Sorter100|16076_ ;
  assign \new_Sorter100|16177_  = \new_Sorter100|16077_  & \new_Sorter100|16078_ ;
  assign \new_Sorter100|16178_  = \new_Sorter100|16077_  | \new_Sorter100|16078_ ;
  assign \new_Sorter100|16179_  = \new_Sorter100|16079_  & \new_Sorter100|16080_ ;
  assign \new_Sorter100|16180_  = \new_Sorter100|16079_  | \new_Sorter100|16080_ ;
  assign \new_Sorter100|16181_  = \new_Sorter100|16081_  & \new_Sorter100|16082_ ;
  assign \new_Sorter100|16182_  = \new_Sorter100|16081_  | \new_Sorter100|16082_ ;
  assign \new_Sorter100|16183_  = \new_Sorter100|16083_  & \new_Sorter100|16084_ ;
  assign \new_Sorter100|16184_  = \new_Sorter100|16083_  | \new_Sorter100|16084_ ;
  assign \new_Sorter100|16185_  = \new_Sorter100|16085_  & \new_Sorter100|16086_ ;
  assign \new_Sorter100|16186_  = \new_Sorter100|16085_  | \new_Sorter100|16086_ ;
  assign \new_Sorter100|16187_  = \new_Sorter100|16087_  & \new_Sorter100|16088_ ;
  assign \new_Sorter100|16188_  = \new_Sorter100|16087_  | \new_Sorter100|16088_ ;
  assign \new_Sorter100|16189_  = \new_Sorter100|16089_  & \new_Sorter100|16090_ ;
  assign \new_Sorter100|16190_  = \new_Sorter100|16089_  | \new_Sorter100|16090_ ;
  assign \new_Sorter100|16191_  = \new_Sorter100|16091_  & \new_Sorter100|16092_ ;
  assign \new_Sorter100|16192_  = \new_Sorter100|16091_  | \new_Sorter100|16092_ ;
  assign \new_Sorter100|16193_  = \new_Sorter100|16093_  & \new_Sorter100|16094_ ;
  assign \new_Sorter100|16194_  = \new_Sorter100|16093_  | \new_Sorter100|16094_ ;
  assign \new_Sorter100|16195_  = \new_Sorter100|16095_  & \new_Sorter100|16096_ ;
  assign \new_Sorter100|16196_  = \new_Sorter100|16095_  | \new_Sorter100|16096_ ;
  assign \new_Sorter100|16197_  = \new_Sorter100|16097_  & \new_Sorter100|16098_ ;
  assign \new_Sorter100|16198_  = \new_Sorter100|16097_  | \new_Sorter100|16098_ ;
  assign \new_Sorter100|16200_  = \new_Sorter100|16100_  & \new_Sorter100|16101_ ;
  assign \new_Sorter100|16201_  = \new_Sorter100|16100_  | \new_Sorter100|16101_ ;
  assign \new_Sorter100|16202_  = \new_Sorter100|16102_  & \new_Sorter100|16103_ ;
  assign \new_Sorter100|16203_  = \new_Sorter100|16102_  | \new_Sorter100|16103_ ;
  assign \new_Sorter100|16204_  = \new_Sorter100|16104_  & \new_Sorter100|16105_ ;
  assign \new_Sorter100|16205_  = \new_Sorter100|16104_  | \new_Sorter100|16105_ ;
  assign \new_Sorter100|16206_  = \new_Sorter100|16106_  & \new_Sorter100|16107_ ;
  assign \new_Sorter100|16207_  = \new_Sorter100|16106_  | \new_Sorter100|16107_ ;
  assign \new_Sorter100|16208_  = \new_Sorter100|16108_  & \new_Sorter100|16109_ ;
  assign \new_Sorter100|16209_  = \new_Sorter100|16108_  | \new_Sorter100|16109_ ;
  assign \new_Sorter100|16210_  = \new_Sorter100|16110_  & \new_Sorter100|16111_ ;
  assign \new_Sorter100|16211_  = \new_Sorter100|16110_  | \new_Sorter100|16111_ ;
  assign \new_Sorter100|16212_  = \new_Sorter100|16112_  & \new_Sorter100|16113_ ;
  assign \new_Sorter100|16213_  = \new_Sorter100|16112_  | \new_Sorter100|16113_ ;
  assign \new_Sorter100|16214_  = \new_Sorter100|16114_  & \new_Sorter100|16115_ ;
  assign \new_Sorter100|16215_  = \new_Sorter100|16114_  | \new_Sorter100|16115_ ;
  assign \new_Sorter100|16216_  = \new_Sorter100|16116_  & \new_Sorter100|16117_ ;
  assign \new_Sorter100|16217_  = \new_Sorter100|16116_  | \new_Sorter100|16117_ ;
  assign \new_Sorter100|16218_  = \new_Sorter100|16118_  & \new_Sorter100|16119_ ;
  assign \new_Sorter100|16219_  = \new_Sorter100|16118_  | \new_Sorter100|16119_ ;
  assign \new_Sorter100|16220_  = \new_Sorter100|16120_  & \new_Sorter100|16121_ ;
  assign \new_Sorter100|16221_  = \new_Sorter100|16120_  | \new_Sorter100|16121_ ;
  assign \new_Sorter100|16222_  = \new_Sorter100|16122_  & \new_Sorter100|16123_ ;
  assign \new_Sorter100|16223_  = \new_Sorter100|16122_  | \new_Sorter100|16123_ ;
  assign \new_Sorter100|16224_  = \new_Sorter100|16124_  & \new_Sorter100|16125_ ;
  assign \new_Sorter100|16225_  = \new_Sorter100|16124_  | \new_Sorter100|16125_ ;
  assign \new_Sorter100|16226_  = \new_Sorter100|16126_  & \new_Sorter100|16127_ ;
  assign \new_Sorter100|16227_  = \new_Sorter100|16126_  | \new_Sorter100|16127_ ;
  assign \new_Sorter100|16228_  = \new_Sorter100|16128_  & \new_Sorter100|16129_ ;
  assign \new_Sorter100|16229_  = \new_Sorter100|16128_  | \new_Sorter100|16129_ ;
  assign \new_Sorter100|16230_  = \new_Sorter100|16130_  & \new_Sorter100|16131_ ;
  assign \new_Sorter100|16231_  = \new_Sorter100|16130_  | \new_Sorter100|16131_ ;
  assign \new_Sorter100|16232_  = \new_Sorter100|16132_  & \new_Sorter100|16133_ ;
  assign \new_Sorter100|16233_  = \new_Sorter100|16132_  | \new_Sorter100|16133_ ;
  assign \new_Sorter100|16234_  = \new_Sorter100|16134_  & \new_Sorter100|16135_ ;
  assign \new_Sorter100|16235_  = \new_Sorter100|16134_  | \new_Sorter100|16135_ ;
  assign \new_Sorter100|16236_  = \new_Sorter100|16136_  & \new_Sorter100|16137_ ;
  assign \new_Sorter100|16237_  = \new_Sorter100|16136_  | \new_Sorter100|16137_ ;
  assign \new_Sorter100|16238_  = \new_Sorter100|16138_  & \new_Sorter100|16139_ ;
  assign \new_Sorter100|16239_  = \new_Sorter100|16138_  | \new_Sorter100|16139_ ;
  assign \new_Sorter100|16240_  = \new_Sorter100|16140_  & \new_Sorter100|16141_ ;
  assign \new_Sorter100|16241_  = \new_Sorter100|16140_  | \new_Sorter100|16141_ ;
  assign \new_Sorter100|16242_  = \new_Sorter100|16142_  & \new_Sorter100|16143_ ;
  assign \new_Sorter100|16243_  = \new_Sorter100|16142_  | \new_Sorter100|16143_ ;
  assign \new_Sorter100|16244_  = \new_Sorter100|16144_  & \new_Sorter100|16145_ ;
  assign \new_Sorter100|16245_  = \new_Sorter100|16144_  | \new_Sorter100|16145_ ;
  assign \new_Sorter100|16246_  = \new_Sorter100|16146_  & \new_Sorter100|16147_ ;
  assign \new_Sorter100|16247_  = \new_Sorter100|16146_  | \new_Sorter100|16147_ ;
  assign \new_Sorter100|16248_  = \new_Sorter100|16148_  & \new_Sorter100|16149_ ;
  assign \new_Sorter100|16249_  = \new_Sorter100|16148_  | \new_Sorter100|16149_ ;
  assign \new_Sorter100|16250_  = \new_Sorter100|16150_  & \new_Sorter100|16151_ ;
  assign \new_Sorter100|16251_  = \new_Sorter100|16150_  | \new_Sorter100|16151_ ;
  assign \new_Sorter100|16252_  = \new_Sorter100|16152_  & \new_Sorter100|16153_ ;
  assign \new_Sorter100|16253_  = \new_Sorter100|16152_  | \new_Sorter100|16153_ ;
  assign \new_Sorter100|16254_  = \new_Sorter100|16154_  & \new_Sorter100|16155_ ;
  assign \new_Sorter100|16255_  = \new_Sorter100|16154_  | \new_Sorter100|16155_ ;
  assign \new_Sorter100|16256_  = \new_Sorter100|16156_  & \new_Sorter100|16157_ ;
  assign \new_Sorter100|16257_  = \new_Sorter100|16156_  | \new_Sorter100|16157_ ;
  assign \new_Sorter100|16258_  = \new_Sorter100|16158_  & \new_Sorter100|16159_ ;
  assign \new_Sorter100|16259_  = \new_Sorter100|16158_  | \new_Sorter100|16159_ ;
  assign \new_Sorter100|16260_  = \new_Sorter100|16160_  & \new_Sorter100|16161_ ;
  assign \new_Sorter100|16261_  = \new_Sorter100|16160_  | \new_Sorter100|16161_ ;
  assign \new_Sorter100|16262_  = \new_Sorter100|16162_  & \new_Sorter100|16163_ ;
  assign \new_Sorter100|16263_  = \new_Sorter100|16162_  | \new_Sorter100|16163_ ;
  assign \new_Sorter100|16264_  = \new_Sorter100|16164_  & \new_Sorter100|16165_ ;
  assign \new_Sorter100|16265_  = \new_Sorter100|16164_  | \new_Sorter100|16165_ ;
  assign \new_Sorter100|16266_  = \new_Sorter100|16166_  & \new_Sorter100|16167_ ;
  assign \new_Sorter100|16267_  = \new_Sorter100|16166_  | \new_Sorter100|16167_ ;
  assign \new_Sorter100|16268_  = \new_Sorter100|16168_  & \new_Sorter100|16169_ ;
  assign \new_Sorter100|16269_  = \new_Sorter100|16168_  | \new_Sorter100|16169_ ;
  assign \new_Sorter100|16270_  = \new_Sorter100|16170_  & \new_Sorter100|16171_ ;
  assign \new_Sorter100|16271_  = \new_Sorter100|16170_  | \new_Sorter100|16171_ ;
  assign \new_Sorter100|16272_  = \new_Sorter100|16172_  & \new_Sorter100|16173_ ;
  assign \new_Sorter100|16273_  = \new_Sorter100|16172_  | \new_Sorter100|16173_ ;
  assign \new_Sorter100|16274_  = \new_Sorter100|16174_  & \new_Sorter100|16175_ ;
  assign \new_Sorter100|16275_  = \new_Sorter100|16174_  | \new_Sorter100|16175_ ;
  assign \new_Sorter100|16276_  = \new_Sorter100|16176_  & \new_Sorter100|16177_ ;
  assign \new_Sorter100|16277_  = \new_Sorter100|16176_  | \new_Sorter100|16177_ ;
  assign \new_Sorter100|16278_  = \new_Sorter100|16178_  & \new_Sorter100|16179_ ;
  assign \new_Sorter100|16279_  = \new_Sorter100|16178_  | \new_Sorter100|16179_ ;
  assign \new_Sorter100|16280_  = \new_Sorter100|16180_  & \new_Sorter100|16181_ ;
  assign \new_Sorter100|16281_  = \new_Sorter100|16180_  | \new_Sorter100|16181_ ;
  assign \new_Sorter100|16282_  = \new_Sorter100|16182_  & \new_Sorter100|16183_ ;
  assign \new_Sorter100|16283_  = \new_Sorter100|16182_  | \new_Sorter100|16183_ ;
  assign \new_Sorter100|16284_  = \new_Sorter100|16184_  & \new_Sorter100|16185_ ;
  assign \new_Sorter100|16285_  = \new_Sorter100|16184_  | \new_Sorter100|16185_ ;
  assign \new_Sorter100|16286_  = \new_Sorter100|16186_  & \new_Sorter100|16187_ ;
  assign \new_Sorter100|16287_  = \new_Sorter100|16186_  | \new_Sorter100|16187_ ;
  assign \new_Sorter100|16288_  = \new_Sorter100|16188_  & \new_Sorter100|16189_ ;
  assign \new_Sorter100|16289_  = \new_Sorter100|16188_  | \new_Sorter100|16189_ ;
  assign \new_Sorter100|16290_  = \new_Sorter100|16190_  & \new_Sorter100|16191_ ;
  assign \new_Sorter100|16291_  = \new_Sorter100|16190_  | \new_Sorter100|16191_ ;
  assign \new_Sorter100|16292_  = \new_Sorter100|16192_  & \new_Sorter100|16193_ ;
  assign \new_Sorter100|16293_  = \new_Sorter100|16192_  | \new_Sorter100|16193_ ;
  assign \new_Sorter100|16294_  = \new_Sorter100|16194_  & \new_Sorter100|16195_ ;
  assign \new_Sorter100|16295_  = \new_Sorter100|16194_  | \new_Sorter100|16195_ ;
  assign \new_Sorter100|16296_  = \new_Sorter100|16196_  & \new_Sorter100|16197_ ;
  assign \new_Sorter100|16297_  = \new_Sorter100|16196_  | \new_Sorter100|16197_ ;
  assign \new_Sorter100|16298_  = \new_Sorter100|16198_  & \new_Sorter100|16199_ ;
  assign \new_Sorter100|16299_  = \new_Sorter100|16198_  | \new_Sorter100|16199_ ;
  assign \new_Sorter100|16300_  = \new_Sorter100|16200_ ;
  assign \new_Sorter100|16399_  = \new_Sorter100|16299_ ;
  assign \new_Sorter100|16301_  = \new_Sorter100|16201_  & \new_Sorter100|16202_ ;
  assign \new_Sorter100|16302_  = \new_Sorter100|16201_  | \new_Sorter100|16202_ ;
  assign \new_Sorter100|16303_  = \new_Sorter100|16203_  & \new_Sorter100|16204_ ;
  assign \new_Sorter100|16304_  = \new_Sorter100|16203_  | \new_Sorter100|16204_ ;
  assign \new_Sorter100|16305_  = \new_Sorter100|16205_  & \new_Sorter100|16206_ ;
  assign \new_Sorter100|16306_  = \new_Sorter100|16205_  | \new_Sorter100|16206_ ;
  assign \new_Sorter100|16307_  = \new_Sorter100|16207_  & \new_Sorter100|16208_ ;
  assign \new_Sorter100|16308_  = \new_Sorter100|16207_  | \new_Sorter100|16208_ ;
  assign \new_Sorter100|16309_  = \new_Sorter100|16209_  & \new_Sorter100|16210_ ;
  assign \new_Sorter100|16310_  = \new_Sorter100|16209_  | \new_Sorter100|16210_ ;
  assign \new_Sorter100|16311_  = \new_Sorter100|16211_  & \new_Sorter100|16212_ ;
  assign \new_Sorter100|16312_  = \new_Sorter100|16211_  | \new_Sorter100|16212_ ;
  assign \new_Sorter100|16313_  = \new_Sorter100|16213_  & \new_Sorter100|16214_ ;
  assign \new_Sorter100|16314_  = \new_Sorter100|16213_  | \new_Sorter100|16214_ ;
  assign \new_Sorter100|16315_  = \new_Sorter100|16215_  & \new_Sorter100|16216_ ;
  assign \new_Sorter100|16316_  = \new_Sorter100|16215_  | \new_Sorter100|16216_ ;
  assign \new_Sorter100|16317_  = \new_Sorter100|16217_  & \new_Sorter100|16218_ ;
  assign \new_Sorter100|16318_  = \new_Sorter100|16217_  | \new_Sorter100|16218_ ;
  assign \new_Sorter100|16319_  = \new_Sorter100|16219_  & \new_Sorter100|16220_ ;
  assign \new_Sorter100|16320_  = \new_Sorter100|16219_  | \new_Sorter100|16220_ ;
  assign \new_Sorter100|16321_  = \new_Sorter100|16221_  & \new_Sorter100|16222_ ;
  assign \new_Sorter100|16322_  = \new_Sorter100|16221_  | \new_Sorter100|16222_ ;
  assign \new_Sorter100|16323_  = \new_Sorter100|16223_  & \new_Sorter100|16224_ ;
  assign \new_Sorter100|16324_  = \new_Sorter100|16223_  | \new_Sorter100|16224_ ;
  assign \new_Sorter100|16325_  = \new_Sorter100|16225_  & \new_Sorter100|16226_ ;
  assign \new_Sorter100|16326_  = \new_Sorter100|16225_  | \new_Sorter100|16226_ ;
  assign \new_Sorter100|16327_  = \new_Sorter100|16227_  & \new_Sorter100|16228_ ;
  assign \new_Sorter100|16328_  = \new_Sorter100|16227_  | \new_Sorter100|16228_ ;
  assign \new_Sorter100|16329_  = \new_Sorter100|16229_  & \new_Sorter100|16230_ ;
  assign \new_Sorter100|16330_  = \new_Sorter100|16229_  | \new_Sorter100|16230_ ;
  assign \new_Sorter100|16331_  = \new_Sorter100|16231_  & \new_Sorter100|16232_ ;
  assign \new_Sorter100|16332_  = \new_Sorter100|16231_  | \new_Sorter100|16232_ ;
  assign \new_Sorter100|16333_  = \new_Sorter100|16233_  & \new_Sorter100|16234_ ;
  assign \new_Sorter100|16334_  = \new_Sorter100|16233_  | \new_Sorter100|16234_ ;
  assign \new_Sorter100|16335_  = \new_Sorter100|16235_  & \new_Sorter100|16236_ ;
  assign \new_Sorter100|16336_  = \new_Sorter100|16235_  | \new_Sorter100|16236_ ;
  assign \new_Sorter100|16337_  = \new_Sorter100|16237_  & \new_Sorter100|16238_ ;
  assign \new_Sorter100|16338_  = \new_Sorter100|16237_  | \new_Sorter100|16238_ ;
  assign \new_Sorter100|16339_  = \new_Sorter100|16239_  & \new_Sorter100|16240_ ;
  assign \new_Sorter100|16340_  = \new_Sorter100|16239_  | \new_Sorter100|16240_ ;
  assign \new_Sorter100|16341_  = \new_Sorter100|16241_  & \new_Sorter100|16242_ ;
  assign \new_Sorter100|16342_  = \new_Sorter100|16241_  | \new_Sorter100|16242_ ;
  assign \new_Sorter100|16343_  = \new_Sorter100|16243_  & \new_Sorter100|16244_ ;
  assign \new_Sorter100|16344_  = \new_Sorter100|16243_  | \new_Sorter100|16244_ ;
  assign \new_Sorter100|16345_  = \new_Sorter100|16245_  & \new_Sorter100|16246_ ;
  assign \new_Sorter100|16346_  = \new_Sorter100|16245_  | \new_Sorter100|16246_ ;
  assign \new_Sorter100|16347_  = \new_Sorter100|16247_  & \new_Sorter100|16248_ ;
  assign \new_Sorter100|16348_  = \new_Sorter100|16247_  | \new_Sorter100|16248_ ;
  assign \new_Sorter100|16349_  = \new_Sorter100|16249_  & \new_Sorter100|16250_ ;
  assign \new_Sorter100|16350_  = \new_Sorter100|16249_  | \new_Sorter100|16250_ ;
  assign \new_Sorter100|16351_  = \new_Sorter100|16251_  & \new_Sorter100|16252_ ;
  assign \new_Sorter100|16352_  = \new_Sorter100|16251_  | \new_Sorter100|16252_ ;
  assign \new_Sorter100|16353_  = \new_Sorter100|16253_  & \new_Sorter100|16254_ ;
  assign \new_Sorter100|16354_  = \new_Sorter100|16253_  | \new_Sorter100|16254_ ;
  assign \new_Sorter100|16355_  = \new_Sorter100|16255_  & \new_Sorter100|16256_ ;
  assign \new_Sorter100|16356_  = \new_Sorter100|16255_  | \new_Sorter100|16256_ ;
  assign \new_Sorter100|16357_  = \new_Sorter100|16257_  & \new_Sorter100|16258_ ;
  assign \new_Sorter100|16358_  = \new_Sorter100|16257_  | \new_Sorter100|16258_ ;
  assign \new_Sorter100|16359_  = \new_Sorter100|16259_  & \new_Sorter100|16260_ ;
  assign \new_Sorter100|16360_  = \new_Sorter100|16259_  | \new_Sorter100|16260_ ;
  assign \new_Sorter100|16361_  = \new_Sorter100|16261_  & \new_Sorter100|16262_ ;
  assign \new_Sorter100|16362_  = \new_Sorter100|16261_  | \new_Sorter100|16262_ ;
  assign \new_Sorter100|16363_  = \new_Sorter100|16263_  & \new_Sorter100|16264_ ;
  assign \new_Sorter100|16364_  = \new_Sorter100|16263_  | \new_Sorter100|16264_ ;
  assign \new_Sorter100|16365_  = \new_Sorter100|16265_  & \new_Sorter100|16266_ ;
  assign \new_Sorter100|16366_  = \new_Sorter100|16265_  | \new_Sorter100|16266_ ;
  assign \new_Sorter100|16367_  = \new_Sorter100|16267_  & \new_Sorter100|16268_ ;
  assign \new_Sorter100|16368_  = \new_Sorter100|16267_  | \new_Sorter100|16268_ ;
  assign \new_Sorter100|16369_  = \new_Sorter100|16269_  & \new_Sorter100|16270_ ;
  assign \new_Sorter100|16370_  = \new_Sorter100|16269_  | \new_Sorter100|16270_ ;
  assign \new_Sorter100|16371_  = \new_Sorter100|16271_  & \new_Sorter100|16272_ ;
  assign \new_Sorter100|16372_  = \new_Sorter100|16271_  | \new_Sorter100|16272_ ;
  assign \new_Sorter100|16373_  = \new_Sorter100|16273_  & \new_Sorter100|16274_ ;
  assign \new_Sorter100|16374_  = \new_Sorter100|16273_  | \new_Sorter100|16274_ ;
  assign \new_Sorter100|16375_  = \new_Sorter100|16275_  & \new_Sorter100|16276_ ;
  assign \new_Sorter100|16376_  = \new_Sorter100|16275_  | \new_Sorter100|16276_ ;
  assign \new_Sorter100|16377_  = \new_Sorter100|16277_  & \new_Sorter100|16278_ ;
  assign \new_Sorter100|16378_  = \new_Sorter100|16277_  | \new_Sorter100|16278_ ;
  assign \new_Sorter100|16379_  = \new_Sorter100|16279_  & \new_Sorter100|16280_ ;
  assign \new_Sorter100|16380_  = \new_Sorter100|16279_  | \new_Sorter100|16280_ ;
  assign \new_Sorter100|16381_  = \new_Sorter100|16281_  & \new_Sorter100|16282_ ;
  assign \new_Sorter100|16382_  = \new_Sorter100|16281_  | \new_Sorter100|16282_ ;
  assign \new_Sorter100|16383_  = \new_Sorter100|16283_  & \new_Sorter100|16284_ ;
  assign \new_Sorter100|16384_  = \new_Sorter100|16283_  | \new_Sorter100|16284_ ;
  assign \new_Sorter100|16385_  = \new_Sorter100|16285_  & \new_Sorter100|16286_ ;
  assign \new_Sorter100|16386_  = \new_Sorter100|16285_  | \new_Sorter100|16286_ ;
  assign \new_Sorter100|16387_  = \new_Sorter100|16287_  & \new_Sorter100|16288_ ;
  assign \new_Sorter100|16388_  = \new_Sorter100|16287_  | \new_Sorter100|16288_ ;
  assign \new_Sorter100|16389_  = \new_Sorter100|16289_  & \new_Sorter100|16290_ ;
  assign \new_Sorter100|16390_  = \new_Sorter100|16289_  | \new_Sorter100|16290_ ;
  assign \new_Sorter100|16391_  = \new_Sorter100|16291_  & \new_Sorter100|16292_ ;
  assign \new_Sorter100|16392_  = \new_Sorter100|16291_  | \new_Sorter100|16292_ ;
  assign \new_Sorter100|16393_  = \new_Sorter100|16293_  & \new_Sorter100|16294_ ;
  assign \new_Sorter100|16394_  = \new_Sorter100|16293_  | \new_Sorter100|16294_ ;
  assign \new_Sorter100|16395_  = \new_Sorter100|16295_  & \new_Sorter100|16296_ ;
  assign \new_Sorter100|16396_  = \new_Sorter100|16295_  | \new_Sorter100|16296_ ;
  assign \new_Sorter100|16397_  = \new_Sorter100|16297_  & \new_Sorter100|16298_ ;
  assign \new_Sorter100|16398_  = \new_Sorter100|16297_  | \new_Sorter100|16298_ ;
  assign \new_Sorter100|16400_  = \new_Sorter100|16300_  & \new_Sorter100|16301_ ;
  assign \new_Sorter100|16401_  = \new_Sorter100|16300_  | \new_Sorter100|16301_ ;
  assign \new_Sorter100|16402_  = \new_Sorter100|16302_  & \new_Sorter100|16303_ ;
  assign \new_Sorter100|16403_  = \new_Sorter100|16302_  | \new_Sorter100|16303_ ;
  assign \new_Sorter100|16404_  = \new_Sorter100|16304_  & \new_Sorter100|16305_ ;
  assign \new_Sorter100|16405_  = \new_Sorter100|16304_  | \new_Sorter100|16305_ ;
  assign \new_Sorter100|16406_  = \new_Sorter100|16306_  & \new_Sorter100|16307_ ;
  assign \new_Sorter100|16407_  = \new_Sorter100|16306_  | \new_Sorter100|16307_ ;
  assign \new_Sorter100|16408_  = \new_Sorter100|16308_  & \new_Sorter100|16309_ ;
  assign \new_Sorter100|16409_  = \new_Sorter100|16308_  | \new_Sorter100|16309_ ;
  assign \new_Sorter100|16410_  = \new_Sorter100|16310_  & \new_Sorter100|16311_ ;
  assign \new_Sorter100|16411_  = \new_Sorter100|16310_  | \new_Sorter100|16311_ ;
  assign \new_Sorter100|16412_  = \new_Sorter100|16312_  & \new_Sorter100|16313_ ;
  assign \new_Sorter100|16413_  = \new_Sorter100|16312_  | \new_Sorter100|16313_ ;
  assign \new_Sorter100|16414_  = \new_Sorter100|16314_  & \new_Sorter100|16315_ ;
  assign \new_Sorter100|16415_  = \new_Sorter100|16314_  | \new_Sorter100|16315_ ;
  assign \new_Sorter100|16416_  = \new_Sorter100|16316_  & \new_Sorter100|16317_ ;
  assign \new_Sorter100|16417_  = \new_Sorter100|16316_  | \new_Sorter100|16317_ ;
  assign \new_Sorter100|16418_  = \new_Sorter100|16318_  & \new_Sorter100|16319_ ;
  assign \new_Sorter100|16419_  = \new_Sorter100|16318_  | \new_Sorter100|16319_ ;
  assign \new_Sorter100|16420_  = \new_Sorter100|16320_  & \new_Sorter100|16321_ ;
  assign \new_Sorter100|16421_  = \new_Sorter100|16320_  | \new_Sorter100|16321_ ;
  assign \new_Sorter100|16422_  = \new_Sorter100|16322_  & \new_Sorter100|16323_ ;
  assign \new_Sorter100|16423_  = \new_Sorter100|16322_  | \new_Sorter100|16323_ ;
  assign \new_Sorter100|16424_  = \new_Sorter100|16324_  & \new_Sorter100|16325_ ;
  assign \new_Sorter100|16425_  = \new_Sorter100|16324_  | \new_Sorter100|16325_ ;
  assign \new_Sorter100|16426_  = \new_Sorter100|16326_  & \new_Sorter100|16327_ ;
  assign \new_Sorter100|16427_  = \new_Sorter100|16326_  | \new_Sorter100|16327_ ;
  assign \new_Sorter100|16428_  = \new_Sorter100|16328_  & \new_Sorter100|16329_ ;
  assign \new_Sorter100|16429_  = \new_Sorter100|16328_  | \new_Sorter100|16329_ ;
  assign \new_Sorter100|16430_  = \new_Sorter100|16330_  & \new_Sorter100|16331_ ;
  assign \new_Sorter100|16431_  = \new_Sorter100|16330_  | \new_Sorter100|16331_ ;
  assign \new_Sorter100|16432_  = \new_Sorter100|16332_  & \new_Sorter100|16333_ ;
  assign \new_Sorter100|16433_  = \new_Sorter100|16332_  | \new_Sorter100|16333_ ;
  assign \new_Sorter100|16434_  = \new_Sorter100|16334_  & \new_Sorter100|16335_ ;
  assign \new_Sorter100|16435_  = \new_Sorter100|16334_  | \new_Sorter100|16335_ ;
  assign \new_Sorter100|16436_  = \new_Sorter100|16336_  & \new_Sorter100|16337_ ;
  assign \new_Sorter100|16437_  = \new_Sorter100|16336_  | \new_Sorter100|16337_ ;
  assign \new_Sorter100|16438_  = \new_Sorter100|16338_  & \new_Sorter100|16339_ ;
  assign \new_Sorter100|16439_  = \new_Sorter100|16338_  | \new_Sorter100|16339_ ;
  assign \new_Sorter100|16440_  = \new_Sorter100|16340_  & \new_Sorter100|16341_ ;
  assign \new_Sorter100|16441_  = \new_Sorter100|16340_  | \new_Sorter100|16341_ ;
  assign \new_Sorter100|16442_  = \new_Sorter100|16342_  & \new_Sorter100|16343_ ;
  assign \new_Sorter100|16443_  = \new_Sorter100|16342_  | \new_Sorter100|16343_ ;
  assign \new_Sorter100|16444_  = \new_Sorter100|16344_  & \new_Sorter100|16345_ ;
  assign \new_Sorter100|16445_  = \new_Sorter100|16344_  | \new_Sorter100|16345_ ;
  assign \new_Sorter100|16446_  = \new_Sorter100|16346_  & \new_Sorter100|16347_ ;
  assign \new_Sorter100|16447_  = \new_Sorter100|16346_  | \new_Sorter100|16347_ ;
  assign \new_Sorter100|16448_  = \new_Sorter100|16348_  & \new_Sorter100|16349_ ;
  assign \new_Sorter100|16449_  = \new_Sorter100|16348_  | \new_Sorter100|16349_ ;
  assign \new_Sorter100|16450_  = \new_Sorter100|16350_  & \new_Sorter100|16351_ ;
  assign \new_Sorter100|16451_  = \new_Sorter100|16350_  | \new_Sorter100|16351_ ;
  assign \new_Sorter100|16452_  = \new_Sorter100|16352_  & \new_Sorter100|16353_ ;
  assign \new_Sorter100|16453_  = \new_Sorter100|16352_  | \new_Sorter100|16353_ ;
  assign \new_Sorter100|16454_  = \new_Sorter100|16354_  & \new_Sorter100|16355_ ;
  assign \new_Sorter100|16455_  = \new_Sorter100|16354_  | \new_Sorter100|16355_ ;
  assign \new_Sorter100|16456_  = \new_Sorter100|16356_  & \new_Sorter100|16357_ ;
  assign \new_Sorter100|16457_  = \new_Sorter100|16356_  | \new_Sorter100|16357_ ;
  assign \new_Sorter100|16458_  = \new_Sorter100|16358_  & \new_Sorter100|16359_ ;
  assign \new_Sorter100|16459_  = \new_Sorter100|16358_  | \new_Sorter100|16359_ ;
  assign \new_Sorter100|16460_  = \new_Sorter100|16360_  & \new_Sorter100|16361_ ;
  assign \new_Sorter100|16461_  = \new_Sorter100|16360_  | \new_Sorter100|16361_ ;
  assign \new_Sorter100|16462_  = \new_Sorter100|16362_  & \new_Sorter100|16363_ ;
  assign \new_Sorter100|16463_  = \new_Sorter100|16362_  | \new_Sorter100|16363_ ;
  assign \new_Sorter100|16464_  = \new_Sorter100|16364_  & \new_Sorter100|16365_ ;
  assign \new_Sorter100|16465_  = \new_Sorter100|16364_  | \new_Sorter100|16365_ ;
  assign \new_Sorter100|16466_  = \new_Sorter100|16366_  & \new_Sorter100|16367_ ;
  assign \new_Sorter100|16467_  = \new_Sorter100|16366_  | \new_Sorter100|16367_ ;
  assign \new_Sorter100|16468_  = \new_Sorter100|16368_  & \new_Sorter100|16369_ ;
  assign \new_Sorter100|16469_  = \new_Sorter100|16368_  | \new_Sorter100|16369_ ;
  assign \new_Sorter100|16470_  = \new_Sorter100|16370_  & \new_Sorter100|16371_ ;
  assign \new_Sorter100|16471_  = \new_Sorter100|16370_  | \new_Sorter100|16371_ ;
  assign \new_Sorter100|16472_  = \new_Sorter100|16372_  & \new_Sorter100|16373_ ;
  assign \new_Sorter100|16473_  = \new_Sorter100|16372_  | \new_Sorter100|16373_ ;
  assign \new_Sorter100|16474_  = \new_Sorter100|16374_  & \new_Sorter100|16375_ ;
  assign \new_Sorter100|16475_  = \new_Sorter100|16374_  | \new_Sorter100|16375_ ;
  assign \new_Sorter100|16476_  = \new_Sorter100|16376_  & \new_Sorter100|16377_ ;
  assign \new_Sorter100|16477_  = \new_Sorter100|16376_  | \new_Sorter100|16377_ ;
  assign \new_Sorter100|16478_  = \new_Sorter100|16378_  & \new_Sorter100|16379_ ;
  assign \new_Sorter100|16479_  = \new_Sorter100|16378_  | \new_Sorter100|16379_ ;
  assign \new_Sorter100|16480_  = \new_Sorter100|16380_  & \new_Sorter100|16381_ ;
  assign \new_Sorter100|16481_  = \new_Sorter100|16380_  | \new_Sorter100|16381_ ;
  assign \new_Sorter100|16482_  = \new_Sorter100|16382_  & \new_Sorter100|16383_ ;
  assign \new_Sorter100|16483_  = \new_Sorter100|16382_  | \new_Sorter100|16383_ ;
  assign \new_Sorter100|16484_  = \new_Sorter100|16384_  & \new_Sorter100|16385_ ;
  assign \new_Sorter100|16485_  = \new_Sorter100|16384_  | \new_Sorter100|16385_ ;
  assign \new_Sorter100|16486_  = \new_Sorter100|16386_  & \new_Sorter100|16387_ ;
  assign \new_Sorter100|16487_  = \new_Sorter100|16386_  | \new_Sorter100|16387_ ;
  assign \new_Sorter100|16488_  = \new_Sorter100|16388_  & \new_Sorter100|16389_ ;
  assign \new_Sorter100|16489_  = \new_Sorter100|16388_  | \new_Sorter100|16389_ ;
  assign \new_Sorter100|16490_  = \new_Sorter100|16390_  & \new_Sorter100|16391_ ;
  assign \new_Sorter100|16491_  = \new_Sorter100|16390_  | \new_Sorter100|16391_ ;
  assign \new_Sorter100|16492_  = \new_Sorter100|16392_  & \new_Sorter100|16393_ ;
  assign \new_Sorter100|16493_  = \new_Sorter100|16392_  | \new_Sorter100|16393_ ;
  assign \new_Sorter100|16494_  = \new_Sorter100|16394_  & \new_Sorter100|16395_ ;
  assign \new_Sorter100|16495_  = \new_Sorter100|16394_  | \new_Sorter100|16395_ ;
  assign \new_Sorter100|16496_  = \new_Sorter100|16396_  & \new_Sorter100|16397_ ;
  assign \new_Sorter100|16497_  = \new_Sorter100|16396_  | \new_Sorter100|16397_ ;
  assign \new_Sorter100|16498_  = \new_Sorter100|16398_  & \new_Sorter100|16399_ ;
  assign \new_Sorter100|16499_  = \new_Sorter100|16398_  | \new_Sorter100|16399_ ;
  assign \new_Sorter100|16500_  = \new_Sorter100|16400_ ;
  assign \new_Sorter100|16599_  = \new_Sorter100|16499_ ;
  assign \new_Sorter100|16501_  = \new_Sorter100|16401_  & \new_Sorter100|16402_ ;
  assign \new_Sorter100|16502_  = \new_Sorter100|16401_  | \new_Sorter100|16402_ ;
  assign \new_Sorter100|16503_  = \new_Sorter100|16403_  & \new_Sorter100|16404_ ;
  assign \new_Sorter100|16504_  = \new_Sorter100|16403_  | \new_Sorter100|16404_ ;
  assign \new_Sorter100|16505_  = \new_Sorter100|16405_  & \new_Sorter100|16406_ ;
  assign \new_Sorter100|16506_  = \new_Sorter100|16405_  | \new_Sorter100|16406_ ;
  assign \new_Sorter100|16507_  = \new_Sorter100|16407_  & \new_Sorter100|16408_ ;
  assign \new_Sorter100|16508_  = \new_Sorter100|16407_  | \new_Sorter100|16408_ ;
  assign \new_Sorter100|16509_  = \new_Sorter100|16409_  & \new_Sorter100|16410_ ;
  assign \new_Sorter100|16510_  = \new_Sorter100|16409_  | \new_Sorter100|16410_ ;
  assign \new_Sorter100|16511_  = \new_Sorter100|16411_  & \new_Sorter100|16412_ ;
  assign \new_Sorter100|16512_  = \new_Sorter100|16411_  | \new_Sorter100|16412_ ;
  assign \new_Sorter100|16513_  = \new_Sorter100|16413_  & \new_Sorter100|16414_ ;
  assign \new_Sorter100|16514_  = \new_Sorter100|16413_  | \new_Sorter100|16414_ ;
  assign \new_Sorter100|16515_  = \new_Sorter100|16415_  & \new_Sorter100|16416_ ;
  assign \new_Sorter100|16516_  = \new_Sorter100|16415_  | \new_Sorter100|16416_ ;
  assign \new_Sorter100|16517_  = \new_Sorter100|16417_  & \new_Sorter100|16418_ ;
  assign \new_Sorter100|16518_  = \new_Sorter100|16417_  | \new_Sorter100|16418_ ;
  assign \new_Sorter100|16519_  = \new_Sorter100|16419_  & \new_Sorter100|16420_ ;
  assign \new_Sorter100|16520_  = \new_Sorter100|16419_  | \new_Sorter100|16420_ ;
  assign \new_Sorter100|16521_  = \new_Sorter100|16421_  & \new_Sorter100|16422_ ;
  assign \new_Sorter100|16522_  = \new_Sorter100|16421_  | \new_Sorter100|16422_ ;
  assign \new_Sorter100|16523_  = \new_Sorter100|16423_  & \new_Sorter100|16424_ ;
  assign \new_Sorter100|16524_  = \new_Sorter100|16423_  | \new_Sorter100|16424_ ;
  assign \new_Sorter100|16525_  = \new_Sorter100|16425_  & \new_Sorter100|16426_ ;
  assign \new_Sorter100|16526_  = \new_Sorter100|16425_  | \new_Sorter100|16426_ ;
  assign \new_Sorter100|16527_  = \new_Sorter100|16427_  & \new_Sorter100|16428_ ;
  assign \new_Sorter100|16528_  = \new_Sorter100|16427_  | \new_Sorter100|16428_ ;
  assign \new_Sorter100|16529_  = \new_Sorter100|16429_  & \new_Sorter100|16430_ ;
  assign \new_Sorter100|16530_  = \new_Sorter100|16429_  | \new_Sorter100|16430_ ;
  assign \new_Sorter100|16531_  = \new_Sorter100|16431_  & \new_Sorter100|16432_ ;
  assign \new_Sorter100|16532_  = \new_Sorter100|16431_  | \new_Sorter100|16432_ ;
  assign \new_Sorter100|16533_  = \new_Sorter100|16433_  & \new_Sorter100|16434_ ;
  assign \new_Sorter100|16534_  = \new_Sorter100|16433_  | \new_Sorter100|16434_ ;
  assign \new_Sorter100|16535_  = \new_Sorter100|16435_  & \new_Sorter100|16436_ ;
  assign \new_Sorter100|16536_  = \new_Sorter100|16435_  | \new_Sorter100|16436_ ;
  assign \new_Sorter100|16537_  = \new_Sorter100|16437_  & \new_Sorter100|16438_ ;
  assign \new_Sorter100|16538_  = \new_Sorter100|16437_  | \new_Sorter100|16438_ ;
  assign \new_Sorter100|16539_  = \new_Sorter100|16439_  & \new_Sorter100|16440_ ;
  assign \new_Sorter100|16540_  = \new_Sorter100|16439_  | \new_Sorter100|16440_ ;
  assign \new_Sorter100|16541_  = \new_Sorter100|16441_  & \new_Sorter100|16442_ ;
  assign \new_Sorter100|16542_  = \new_Sorter100|16441_  | \new_Sorter100|16442_ ;
  assign \new_Sorter100|16543_  = \new_Sorter100|16443_  & \new_Sorter100|16444_ ;
  assign \new_Sorter100|16544_  = \new_Sorter100|16443_  | \new_Sorter100|16444_ ;
  assign \new_Sorter100|16545_  = \new_Sorter100|16445_  & \new_Sorter100|16446_ ;
  assign \new_Sorter100|16546_  = \new_Sorter100|16445_  | \new_Sorter100|16446_ ;
  assign \new_Sorter100|16547_  = \new_Sorter100|16447_  & \new_Sorter100|16448_ ;
  assign \new_Sorter100|16548_  = \new_Sorter100|16447_  | \new_Sorter100|16448_ ;
  assign \new_Sorter100|16549_  = \new_Sorter100|16449_  & \new_Sorter100|16450_ ;
  assign \new_Sorter100|16550_  = \new_Sorter100|16449_  | \new_Sorter100|16450_ ;
  assign \new_Sorter100|16551_  = \new_Sorter100|16451_  & \new_Sorter100|16452_ ;
  assign \new_Sorter100|16552_  = \new_Sorter100|16451_  | \new_Sorter100|16452_ ;
  assign \new_Sorter100|16553_  = \new_Sorter100|16453_  & \new_Sorter100|16454_ ;
  assign \new_Sorter100|16554_  = \new_Sorter100|16453_  | \new_Sorter100|16454_ ;
  assign \new_Sorter100|16555_  = \new_Sorter100|16455_  & \new_Sorter100|16456_ ;
  assign \new_Sorter100|16556_  = \new_Sorter100|16455_  | \new_Sorter100|16456_ ;
  assign \new_Sorter100|16557_  = \new_Sorter100|16457_  & \new_Sorter100|16458_ ;
  assign \new_Sorter100|16558_  = \new_Sorter100|16457_  | \new_Sorter100|16458_ ;
  assign \new_Sorter100|16559_  = \new_Sorter100|16459_  & \new_Sorter100|16460_ ;
  assign \new_Sorter100|16560_  = \new_Sorter100|16459_  | \new_Sorter100|16460_ ;
  assign \new_Sorter100|16561_  = \new_Sorter100|16461_  & \new_Sorter100|16462_ ;
  assign \new_Sorter100|16562_  = \new_Sorter100|16461_  | \new_Sorter100|16462_ ;
  assign \new_Sorter100|16563_  = \new_Sorter100|16463_  & \new_Sorter100|16464_ ;
  assign \new_Sorter100|16564_  = \new_Sorter100|16463_  | \new_Sorter100|16464_ ;
  assign \new_Sorter100|16565_  = \new_Sorter100|16465_  & \new_Sorter100|16466_ ;
  assign \new_Sorter100|16566_  = \new_Sorter100|16465_  | \new_Sorter100|16466_ ;
  assign \new_Sorter100|16567_  = \new_Sorter100|16467_  & \new_Sorter100|16468_ ;
  assign \new_Sorter100|16568_  = \new_Sorter100|16467_  | \new_Sorter100|16468_ ;
  assign \new_Sorter100|16569_  = \new_Sorter100|16469_  & \new_Sorter100|16470_ ;
  assign \new_Sorter100|16570_  = \new_Sorter100|16469_  | \new_Sorter100|16470_ ;
  assign \new_Sorter100|16571_  = \new_Sorter100|16471_  & \new_Sorter100|16472_ ;
  assign \new_Sorter100|16572_  = \new_Sorter100|16471_  | \new_Sorter100|16472_ ;
  assign \new_Sorter100|16573_  = \new_Sorter100|16473_  & \new_Sorter100|16474_ ;
  assign \new_Sorter100|16574_  = \new_Sorter100|16473_  | \new_Sorter100|16474_ ;
  assign \new_Sorter100|16575_  = \new_Sorter100|16475_  & \new_Sorter100|16476_ ;
  assign \new_Sorter100|16576_  = \new_Sorter100|16475_  | \new_Sorter100|16476_ ;
  assign \new_Sorter100|16577_  = \new_Sorter100|16477_  & \new_Sorter100|16478_ ;
  assign \new_Sorter100|16578_  = \new_Sorter100|16477_  | \new_Sorter100|16478_ ;
  assign \new_Sorter100|16579_  = \new_Sorter100|16479_  & \new_Sorter100|16480_ ;
  assign \new_Sorter100|16580_  = \new_Sorter100|16479_  | \new_Sorter100|16480_ ;
  assign \new_Sorter100|16581_  = \new_Sorter100|16481_  & \new_Sorter100|16482_ ;
  assign \new_Sorter100|16582_  = \new_Sorter100|16481_  | \new_Sorter100|16482_ ;
  assign \new_Sorter100|16583_  = \new_Sorter100|16483_  & \new_Sorter100|16484_ ;
  assign \new_Sorter100|16584_  = \new_Sorter100|16483_  | \new_Sorter100|16484_ ;
  assign \new_Sorter100|16585_  = \new_Sorter100|16485_  & \new_Sorter100|16486_ ;
  assign \new_Sorter100|16586_  = \new_Sorter100|16485_  | \new_Sorter100|16486_ ;
  assign \new_Sorter100|16587_  = \new_Sorter100|16487_  & \new_Sorter100|16488_ ;
  assign \new_Sorter100|16588_  = \new_Sorter100|16487_  | \new_Sorter100|16488_ ;
  assign \new_Sorter100|16589_  = \new_Sorter100|16489_  & \new_Sorter100|16490_ ;
  assign \new_Sorter100|16590_  = \new_Sorter100|16489_  | \new_Sorter100|16490_ ;
  assign \new_Sorter100|16591_  = \new_Sorter100|16491_  & \new_Sorter100|16492_ ;
  assign \new_Sorter100|16592_  = \new_Sorter100|16491_  | \new_Sorter100|16492_ ;
  assign \new_Sorter100|16593_  = \new_Sorter100|16493_  & \new_Sorter100|16494_ ;
  assign \new_Sorter100|16594_  = \new_Sorter100|16493_  | \new_Sorter100|16494_ ;
  assign \new_Sorter100|16595_  = \new_Sorter100|16495_  & \new_Sorter100|16496_ ;
  assign \new_Sorter100|16596_  = \new_Sorter100|16495_  | \new_Sorter100|16496_ ;
  assign \new_Sorter100|16597_  = \new_Sorter100|16497_  & \new_Sorter100|16498_ ;
  assign \new_Sorter100|16598_  = \new_Sorter100|16497_  | \new_Sorter100|16498_ ;
  assign \new_Sorter100|16600_  = \new_Sorter100|16500_  & \new_Sorter100|16501_ ;
  assign \new_Sorter100|16601_  = \new_Sorter100|16500_  | \new_Sorter100|16501_ ;
  assign \new_Sorter100|16602_  = \new_Sorter100|16502_  & \new_Sorter100|16503_ ;
  assign \new_Sorter100|16603_  = \new_Sorter100|16502_  | \new_Sorter100|16503_ ;
  assign \new_Sorter100|16604_  = \new_Sorter100|16504_  & \new_Sorter100|16505_ ;
  assign \new_Sorter100|16605_  = \new_Sorter100|16504_  | \new_Sorter100|16505_ ;
  assign \new_Sorter100|16606_  = \new_Sorter100|16506_  & \new_Sorter100|16507_ ;
  assign \new_Sorter100|16607_  = \new_Sorter100|16506_  | \new_Sorter100|16507_ ;
  assign \new_Sorter100|16608_  = \new_Sorter100|16508_  & \new_Sorter100|16509_ ;
  assign \new_Sorter100|16609_  = \new_Sorter100|16508_  | \new_Sorter100|16509_ ;
  assign \new_Sorter100|16610_  = \new_Sorter100|16510_  & \new_Sorter100|16511_ ;
  assign \new_Sorter100|16611_  = \new_Sorter100|16510_  | \new_Sorter100|16511_ ;
  assign \new_Sorter100|16612_  = \new_Sorter100|16512_  & \new_Sorter100|16513_ ;
  assign \new_Sorter100|16613_  = \new_Sorter100|16512_  | \new_Sorter100|16513_ ;
  assign \new_Sorter100|16614_  = \new_Sorter100|16514_  & \new_Sorter100|16515_ ;
  assign \new_Sorter100|16615_  = \new_Sorter100|16514_  | \new_Sorter100|16515_ ;
  assign \new_Sorter100|16616_  = \new_Sorter100|16516_  & \new_Sorter100|16517_ ;
  assign \new_Sorter100|16617_  = \new_Sorter100|16516_  | \new_Sorter100|16517_ ;
  assign \new_Sorter100|16618_  = \new_Sorter100|16518_  & \new_Sorter100|16519_ ;
  assign \new_Sorter100|16619_  = \new_Sorter100|16518_  | \new_Sorter100|16519_ ;
  assign \new_Sorter100|16620_  = \new_Sorter100|16520_  & \new_Sorter100|16521_ ;
  assign \new_Sorter100|16621_  = \new_Sorter100|16520_  | \new_Sorter100|16521_ ;
  assign \new_Sorter100|16622_  = \new_Sorter100|16522_  & \new_Sorter100|16523_ ;
  assign \new_Sorter100|16623_  = \new_Sorter100|16522_  | \new_Sorter100|16523_ ;
  assign \new_Sorter100|16624_  = \new_Sorter100|16524_  & \new_Sorter100|16525_ ;
  assign \new_Sorter100|16625_  = \new_Sorter100|16524_  | \new_Sorter100|16525_ ;
  assign \new_Sorter100|16626_  = \new_Sorter100|16526_  & \new_Sorter100|16527_ ;
  assign \new_Sorter100|16627_  = \new_Sorter100|16526_  | \new_Sorter100|16527_ ;
  assign \new_Sorter100|16628_  = \new_Sorter100|16528_  & \new_Sorter100|16529_ ;
  assign \new_Sorter100|16629_  = \new_Sorter100|16528_  | \new_Sorter100|16529_ ;
  assign \new_Sorter100|16630_  = \new_Sorter100|16530_  & \new_Sorter100|16531_ ;
  assign \new_Sorter100|16631_  = \new_Sorter100|16530_  | \new_Sorter100|16531_ ;
  assign \new_Sorter100|16632_  = \new_Sorter100|16532_  & \new_Sorter100|16533_ ;
  assign \new_Sorter100|16633_  = \new_Sorter100|16532_  | \new_Sorter100|16533_ ;
  assign \new_Sorter100|16634_  = \new_Sorter100|16534_  & \new_Sorter100|16535_ ;
  assign \new_Sorter100|16635_  = \new_Sorter100|16534_  | \new_Sorter100|16535_ ;
  assign \new_Sorter100|16636_  = \new_Sorter100|16536_  & \new_Sorter100|16537_ ;
  assign \new_Sorter100|16637_  = \new_Sorter100|16536_  | \new_Sorter100|16537_ ;
  assign \new_Sorter100|16638_  = \new_Sorter100|16538_  & \new_Sorter100|16539_ ;
  assign \new_Sorter100|16639_  = \new_Sorter100|16538_  | \new_Sorter100|16539_ ;
  assign \new_Sorter100|16640_  = \new_Sorter100|16540_  & \new_Sorter100|16541_ ;
  assign \new_Sorter100|16641_  = \new_Sorter100|16540_  | \new_Sorter100|16541_ ;
  assign \new_Sorter100|16642_  = \new_Sorter100|16542_  & \new_Sorter100|16543_ ;
  assign \new_Sorter100|16643_  = \new_Sorter100|16542_  | \new_Sorter100|16543_ ;
  assign \new_Sorter100|16644_  = \new_Sorter100|16544_  & \new_Sorter100|16545_ ;
  assign \new_Sorter100|16645_  = \new_Sorter100|16544_  | \new_Sorter100|16545_ ;
  assign \new_Sorter100|16646_  = \new_Sorter100|16546_  & \new_Sorter100|16547_ ;
  assign \new_Sorter100|16647_  = \new_Sorter100|16546_  | \new_Sorter100|16547_ ;
  assign \new_Sorter100|16648_  = \new_Sorter100|16548_  & \new_Sorter100|16549_ ;
  assign \new_Sorter100|16649_  = \new_Sorter100|16548_  | \new_Sorter100|16549_ ;
  assign \new_Sorter100|16650_  = \new_Sorter100|16550_  & \new_Sorter100|16551_ ;
  assign \new_Sorter100|16651_  = \new_Sorter100|16550_  | \new_Sorter100|16551_ ;
  assign \new_Sorter100|16652_  = \new_Sorter100|16552_  & \new_Sorter100|16553_ ;
  assign \new_Sorter100|16653_  = \new_Sorter100|16552_  | \new_Sorter100|16553_ ;
  assign \new_Sorter100|16654_  = \new_Sorter100|16554_  & \new_Sorter100|16555_ ;
  assign \new_Sorter100|16655_  = \new_Sorter100|16554_  | \new_Sorter100|16555_ ;
  assign \new_Sorter100|16656_  = \new_Sorter100|16556_  & \new_Sorter100|16557_ ;
  assign \new_Sorter100|16657_  = \new_Sorter100|16556_  | \new_Sorter100|16557_ ;
  assign \new_Sorter100|16658_  = \new_Sorter100|16558_  & \new_Sorter100|16559_ ;
  assign \new_Sorter100|16659_  = \new_Sorter100|16558_  | \new_Sorter100|16559_ ;
  assign \new_Sorter100|16660_  = \new_Sorter100|16560_  & \new_Sorter100|16561_ ;
  assign \new_Sorter100|16661_  = \new_Sorter100|16560_  | \new_Sorter100|16561_ ;
  assign \new_Sorter100|16662_  = \new_Sorter100|16562_  & \new_Sorter100|16563_ ;
  assign \new_Sorter100|16663_  = \new_Sorter100|16562_  | \new_Sorter100|16563_ ;
  assign \new_Sorter100|16664_  = \new_Sorter100|16564_  & \new_Sorter100|16565_ ;
  assign \new_Sorter100|16665_  = \new_Sorter100|16564_  | \new_Sorter100|16565_ ;
  assign \new_Sorter100|16666_  = \new_Sorter100|16566_  & \new_Sorter100|16567_ ;
  assign \new_Sorter100|16667_  = \new_Sorter100|16566_  | \new_Sorter100|16567_ ;
  assign \new_Sorter100|16668_  = \new_Sorter100|16568_  & \new_Sorter100|16569_ ;
  assign \new_Sorter100|16669_  = \new_Sorter100|16568_  | \new_Sorter100|16569_ ;
  assign \new_Sorter100|16670_  = \new_Sorter100|16570_  & \new_Sorter100|16571_ ;
  assign \new_Sorter100|16671_  = \new_Sorter100|16570_  | \new_Sorter100|16571_ ;
  assign \new_Sorter100|16672_  = \new_Sorter100|16572_  & \new_Sorter100|16573_ ;
  assign \new_Sorter100|16673_  = \new_Sorter100|16572_  | \new_Sorter100|16573_ ;
  assign \new_Sorter100|16674_  = \new_Sorter100|16574_  & \new_Sorter100|16575_ ;
  assign \new_Sorter100|16675_  = \new_Sorter100|16574_  | \new_Sorter100|16575_ ;
  assign \new_Sorter100|16676_  = \new_Sorter100|16576_  & \new_Sorter100|16577_ ;
  assign \new_Sorter100|16677_  = \new_Sorter100|16576_  | \new_Sorter100|16577_ ;
  assign \new_Sorter100|16678_  = \new_Sorter100|16578_  & \new_Sorter100|16579_ ;
  assign \new_Sorter100|16679_  = \new_Sorter100|16578_  | \new_Sorter100|16579_ ;
  assign \new_Sorter100|16680_  = \new_Sorter100|16580_  & \new_Sorter100|16581_ ;
  assign \new_Sorter100|16681_  = \new_Sorter100|16580_  | \new_Sorter100|16581_ ;
  assign \new_Sorter100|16682_  = \new_Sorter100|16582_  & \new_Sorter100|16583_ ;
  assign \new_Sorter100|16683_  = \new_Sorter100|16582_  | \new_Sorter100|16583_ ;
  assign \new_Sorter100|16684_  = \new_Sorter100|16584_  & \new_Sorter100|16585_ ;
  assign \new_Sorter100|16685_  = \new_Sorter100|16584_  | \new_Sorter100|16585_ ;
  assign \new_Sorter100|16686_  = \new_Sorter100|16586_  & \new_Sorter100|16587_ ;
  assign \new_Sorter100|16687_  = \new_Sorter100|16586_  | \new_Sorter100|16587_ ;
  assign \new_Sorter100|16688_  = \new_Sorter100|16588_  & \new_Sorter100|16589_ ;
  assign \new_Sorter100|16689_  = \new_Sorter100|16588_  | \new_Sorter100|16589_ ;
  assign \new_Sorter100|16690_  = \new_Sorter100|16590_  & \new_Sorter100|16591_ ;
  assign \new_Sorter100|16691_  = \new_Sorter100|16590_  | \new_Sorter100|16591_ ;
  assign \new_Sorter100|16692_  = \new_Sorter100|16592_  & \new_Sorter100|16593_ ;
  assign \new_Sorter100|16693_  = \new_Sorter100|16592_  | \new_Sorter100|16593_ ;
  assign \new_Sorter100|16694_  = \new_Sorter100|16594_  & \new_Sorter100|16595_ ;
  assign \new_Sorter100|16695_  = \new_Sorter100|16594_  | \new_Sorter100|16595_ ;
  assign \new_Sorter100|16696_  = \new_Sorter100|16596_  & \new_Sorter100|16597_ ;
  assign \new_Sorter100|16697_  = \new_Sorter100|16596_  | \new_Sorter100|16597_ ;
  assign \new_Sorter100|16698_  = \new_Sorter100|16598_  & \new_Sorter100|16599_ ;
  assign \new_Sorter100|16699_  = \new_Sorter100|16598_  | \new_Sorter100|16599_ ;
  assign \new_Sorter100|16700_  = \new_Sorter100|16600_ ;
  assign \new_Sorter100|16799_  = \new_Sorter100|16699_ ;
  assign \new_Sorter100|16701_  = \new_Sorter100|16601_  & \new_Sorter100|16602_ ;
  assign \new_Sorter100|16702_  = \new_Sorter100|16601_  | \new_Sorter100|16602_ ;
  assign \new_Sorter100|16703_  = \new_Sorter100|16603_  & \new_Sorter100|16604_ ;
  assign \new_Sorter100|16704_  = \new_Sorter100|16603_  | \new_Sorter100|16604_ ;
  assign \new_Sorter100|16705_  = \new_Sorter100|16605_  & \new_Sorter100|16606_ ;
  assign \new_Sorter100|16706_  = \new_Sorter100|16605_  | \new_Sorter100|16606_ ;
  assign \new_Sorter100|16707_  = \new_Sorter100|16607_  & \new_Sorter100|16608_ ;
  assign \new_Sorter100|16708_  = \new_Sorter100|16607_  | \new_Sorter100|16608_ ;
  assign \new_Sorter100|16709_  = \new_Sorter100|16609_  & \new_Sorter100|16610_ ;
  assign \new_Sorter100|16710_  = \new_Sorter100|16609_  | \new_Sorter100|16610_ ;
  assign \new_Sorter100|16711_  = \new_Sorter100|16611_  & \new_Sorter100|16612_ ;
  assign \new_Sorter100|16712_  = \new_Sorter100|16611_  | \new_Sorter100|16612_ ;
  assign \new_Sorter100|16713_  = \new_Sorter100|16613_  & \new_Sorter100|16614_ ;
  assign \new_Sorter100|16714_  = \new_Sorter100|16613_  | \new_Sorter100|16614_ ;
  assign \new_Sorter100|16715_  = \new_Sorter100|16615_  & \new_Sorter100|16616_ ;
  assign \new_Sorter100|16716_  = \new_Sorter100|16615_  | \new_Sorter100|16616_ ;
  assign \new_Sorter100|16717_  = \new_Sorter100|16617_  & \new_Sorter100|16618_ ;
  assign \new_Sorter100|16718_  = \new_Sorter100|16617_  | \new_Sorter100|16618_ ;
  assign \new_Sorter100|16719_  = \new_Sorter100|16619_  & \new_Sorter100|16620_ ;
  assign \new_Sorter100|16720_  = \new_Sorter100|16619_  | \new_Sorter100|16620_ ;
  assign \new_Sorter100|16721_  = \new_Sorter100|16621_  & \new_Sorter100|16622_ ;
  assign \new_Sorter100|16722_  = \new_Sorter100|16621_  | \new_Sorter100|16622_ ;
  assign \new_Sorter100|16723_  = \new_Sorter100|16623_  & \new_Sorter100|16624_ ;
  assign \new_Sorter100|16724_  = \new_Sorter100|16623_  | \new_Sorter100|16624_ ;
  assign \new_Sorter100|16725_  = \new_Sorter100|16625_  & \new_Sorter100|16626_ ;
  assign \new_Sorter100|16726_  = \new_Sorter100|16625_  | \new_Sorter100|16626_ ;
  assign \new_Sorter100|16727_  = \new_Sorter100|16627_  & \new_Sorter100|16628_ ;
  assign \new_Sorter100|16728_  = \new_Sorter100|16627_  | \new_Sorter100|16628_ ;
  assign \new_Sorter100|16729_  = \new_Sorter100|16629_  & \new_Sorter100|16630_ ;
  assign \new_Sorter100|16730_  = \new_Sorter100|16629_  | \new_Sorter100|16630_ ;
  assign \new_Sorter100|16731_  = \new_Sorter100|16631_  & \new_Sorter100|16632_ ;
  assign \new_Sorter100|16732_  = \new_Sorter100|16631_  | \new_Sorter100|16632_ ;
  assign \new_Sorter100|16733_  = \new_Sorter100|16633_  & \new_Sorter100|16634_ ;
  assign \new_Sorter100|16734_  = \new_Sorter100|16633_  | \new_Sorter100|16634_ ;
  assign \new_Sorter100|16735_  = \new_Sorter100|16635_  & \new_Sorter100|16636_ ;
  assign \new_Sorter100|16736_  = \new_Sorter100|16635_  | \new_Sorter100|16636_ ;
  assign \new_Sorter100|16737_  = \new_Sorter100|16637_  & \new_Sorter100|16638_ ;
  assign \new_Sorter100|16738_  = \new_Sorter100|16637_  | \new_Sorter100|16638_ ;
  assign \new_Sorter100|16739_  = \new_Sorter100|16639_  & \new_Sorter100|16640_ ;
  assign \new_Sorter100|16740_  = \new_Sorter100|16639_  | \new_Sorter100|16640_ ;
  assign \new_Sorter100|16741_  = \new_Sorter100|16641_  & \new_Sorter100|16642_ ;
  assign \new_Sorter100|16742_  = \new_Sorter100|16641_  | \new_Sorter100|16642_ ;
  assign \new_Sorter100|16743_  = \new_Sorter100|16643_  & \new_Sorter100|16644_ ;
  assign \new_Sorter100|16744_  = \new_Sorter100|16643_  | \new_Sorter100|16644_ ;
  assign \new_Sorter100|16745_  = \new_Sorter100|16645_  & \new_Sorter100|16646_ ;
  assign \new_Sorter100|16746_  = \new_Sorter100|16645_  | \new_Sorter100|16646_ ;
  assign \new_Sorter100|16747_  = \new_Sorter100|16647_  & \new_Sorter100|16648_ ;
  assign \new_Sorter100|16748_  = \new_Sorter100|16647_  | \new_Sorter100|16648_ ;
  assign \new_Sorter100|16749_  = \new_Sorter100|16649_  & \new_Sorter100|16650_ ;
  assign \new_Sorter100|16750_  = \new_Sorter100|16649_  | \new_Sorter100|16650_ ;
  assign \new_Sorter100|16751_  = \new_Sorter100|16651_  & \new_Sorter100|16652_ ;
  assign \new_Sorter100|16752_  = \new_Sorter100|16651_  | \new_Sorter100|16652_ ;
  assign \new_Sorter100|16753_  = \new_Sorter100|16653_  & \new_Sorter100|16654_ ;
  assign \new_Sorter100|16754_  = \new_Sorter100|16653_  | \new_Sorter100|16654_ ;
  assign \new_Sorter100|16755_  = \new_Sorter100|16655_  & \new_Sorter100|16656_ ;
  assign \new_Sorter100|16756_  = \new_Sorter100|16655_  | \new_Sorter100|16656_ ;
  assign \new_Sorter100|16757_  = \new_Sorter100|16657_  & \new_Sorter100|16658_ ;
  assign \new_Sorter100|16758_  = \new_Sorter100|16657_  | \new_Sorter100|16658_ ;
  assign \new_Sorter100|16759_  = \new_Sorter100|16659_  & \new_Sorter100|16660_ ;
  assign \new_Sorter100|16760_  = \new_Sorter100|16659_  | \new_Sorter100|16660_ ;
  assign \new_Sorter100|16761_  = \new_Sorter100|16661_  & \new_Sorter100|16662_ ;
  assign \new_Sorter100|16762_  = \new_Sorter100|16661_  | \new_Sorter100|16662_ ;
  assign \new_Sorter100|16763_  = \new_Sorter100|16663_  & \new_Sorter100|16664_ ;
  assign \new_Sorter100|16764_  = \new_Sorter100|16663_  | \new_Sorter100|16664_ ;
  assign \new_Sorter100|16765_  = \new_Sorter100|16665_  & \new_Sorter100|16666_ ;
  assign \new_Sorter100|16766_  = \new_Sorter100|16665_  | \new_Sorter100|16666_ ;
  assign \new_Sorter100|16767_  = \new_Sorter100|16667_  & \new_Sorter100|16668_ ;
  assign \new_Sorter100|16768_  = \new_Sorter100|16667_  | \new_Sorter100|16668_ ;
  assign \new_Sorter100|16769_  = \new_Sorter100|16669_  & \new_Sorter100|16670_ ;
  assign \new_Sorter100|16770_  = \new_Sorter100|16669_  | \new_Sorter100|16670_ ;
  assign \new_Sorter100|16771_  = \new_Sorter100|16671_  & \new_Sorter100|16672_ ;
  assign \new_Sorter100|16772_  = \new_Sorter100|16671_  | \new_Sorter100|16672_ ;
  assign \new_Sorter100|16773_  = \new_Sorter100|16673_  & \new_Sorter100|16674_ ;
  assign \new_Sorter100|16774_  = \new_Sorter100|16673_  | \new_Sorter100|16674_ ;
  assign \new_Sorter100|16775_  = \new_Sorter100|16675_  & \new_Sorter100|16676_ ;
  assign \new_Sorter100|16776_  = \new_Sorter100|16675_  | \new_Sorter100|16676_ ;
  assign \new_Sorter100|16777_  = \new_Sorter100|16677_  & \new_Sorter100|16678_ ;
  assign \new_Sorter100|16778_  = \new_Sorter100|16677_  | \new_Sorter100|16678_ ;
  assign \new_Sorter100|16779_  = \new_Sorter100|16679_  & \new_Sorter100|16680_ ;
  assign \new_Sorter100|16780_  = \new_Sorter100|16679_  | \new_Sorter100|16680_ ;
  assign \new_Sorter100|16781_  = \new_Sorter100|16681_  & \new_Sorter100|16682_ ;
  assign \new_Sorter100|16782_  = \new_Sorter100|16681_  | \new_Sorter100|16682_ ;
  assign \new_Sorter100|16783_  = \new_Sorter100|16683_  & \new_Sorter100|16684_ ;
  assign \new_Sorter100|16784_  = \new_Sorter100|16683_  | \new_Sorter100|16684_ ;
  assign \new_Sorter100|16785_  = \new_Sorter100|16685_  & \new_Sorter100|16686_ ;
  assign \new_Sorter100|16786_  = \new_Sorter100|16685_  | \new_Sorter100|16686_ ;
  assign \new_Sorter100|16787_  = \new_Sorter100|16687_  & \new_Sorter100|16688_ ;
  assign \new_Sorter100|16788_  = \new_Sorter100|16687_  | \new_Sorter100|16688_ ;
  assign \new_Sorter100|16789_  = \new_Sorter100|16689_  & \new_Sorter100|16690_ ;
  assign \new_Sorter100|16790_  = \new_Sorter100|16689_  | \new_Sorter100|16690_ ;
  assign \new_Sorter100|16791_  = \new_Sorter100|16691_  & \new_Sorter100|16692_ ;
  assign \new_Sorter100|16792_  = \new_Sorter100|16691_  | \new_Sorter100|16692_ ;
  assign \new_Sorter100|16793_  = \new_Sorter100|16693_  & \new_Sorter100|16694_ ;
  assign \new_Sorter100|16794_  = \new_Sorter100|16693_  | \new_Sorter100|16694_ ;
  assign \new_Sorter100|16795_  = \new_Sorter100|16695_  & \new_Sorter100|16696_ ;
  assign \new_Sorter100|16796_  = \new_Sorter100|16695_  | \new_Sorter100|16696_ ;
  assign \new_Sorter100|16797_  = \new_Sorter100|16697_  & \new_Sorter100|16698_ ;
  assign \new_Sorter100|16798_  = \new_Sorter100|16697_  | \new_Sorter100|16698_ ;
  assign \new_Sorter100|16800_  = \new_Sorter100|16700_  & \new_Sorter100|16701_ ;
  assign \new_Sorter100|16801_  = \new_Sorter100|16700_  | \new_Sorter100|16701_ ;
  assign \new_Sorter100|16802_  = \new_Sorter100|16702_  & \new_Sorter100|16703_ ;
  assign \new_Sorter100|16803_  = \new_Sorter100|16702_  | \new_Sorter100|16703_ ;
  assign \new_Sorter100|16804_  = \new_Sorter100|16704_  & \new_Sorter100|16705_ ;
  assign \new_Sorter100|16805_  = \new_Sorter100|16704_  | \new_Sorter100|16705_ ;
  assign \new_Sorter100|16806_  = \new_Sorter100|16706_  & \new_Sorter100|16707_ ;
  assign \new_Sorter100|16807_  = \new_Sorter100|16706_  | \new_Sorter100|16707_ ;
  assign \new_Sorter100|16808_  = \new_Sorter100|16708_  & \new_Sorter100|16709_ ;
  assign \new_Sorter100|16809_  = \new_Sorter100|16708_  | \new_Sorter100|16709_ ;
  assign \new_Sorter100|16810_  = \new_Sorter100|16710_  & \new_Sorter100|16711_ ;
  assign \new_Sorter100|16811_  = \new_Sorter100|16710_  | \new_Sorter100|16711_ ;
  assign \new_Sorter100|16812_  = \new_Sorter100|16712_  & \new_Sorter100|16713_ ;
  assign \new_Sorter100|16813_  = \new_Sorter100|16712_  | \new_Sorter100|16713_ ;
  assign \new_Sorter100|16814_  = \new_Sorter100|16714_  & \new_Sorter100|16715_ ;
  assign \new_Sorter100|16815_  = \new_Sorter100|16714_  | \new_Sorter100|16715_ ;
  assign \new_Sorter100|16816_  = \new_Sorter100|16716_  & \new_Sorter100|16717_ ;
  assign \new_Sorter100|16817_  = \new_Sorter100|16716_  | \new_Sorter100|16717_ ;
  assign \new_Sorter100|16818_  = \new_Sorter100|16718_  & \new_Sorter100|16719_ ;
  assign \new_Sorter100|16819_  = \new_Sorter100|16718_  | \new_Sorter100|16719_ ;
  assign \new_Sorter100|16820_  = \new_Sorter100|16720_  & \new_Sorter100|16721_ ;
  assign \new_Sorter100|16821_  = \new_Sorter100|16720_  | \new_Sorter100|16721_ ;
  assign \new_Sorter100|16822_  = \new_Sorter100|16722_  & \new_Sorter100|16723_ ;
  assign \new_Sorter100|16823_  = \new_Sorter100|16722_  | \new_Sorter100|16723_ ;
  assign \new_Sorter100|16824_  = \new_Sorter100|16724_  & \new_Sorter100|16725_ ;
  assign \new_Sorter100|16825_  = \new_Sorter100|16724_  | \new_Sorter100|16725_ ;
  assign \new_Sorter100|16826_  = \new_Sorter100|16726_  & \new_Sorter100|16727_ ;
  assign \new_Sorter100|16827_  = \new_Sorter100|16726_  | \new_Sorter100|16727_ ;
  assign \new_Sorter100|16828_  = \new_Sorter100|16728_  & \new_Sorter100|16729_ ;
  assign \new_Sorter100|16829_  = \new_Sorter100|16728_  | \new_Sorter100|16729_ ;
  assign \new_Sorter100|16830_  = \new_Sorter100|16730_  & \new_Sorter100|16731_ ;
  assign \new_Sorter100|16831_  = \new_Sorter100|16730_  | \new_Sorter100|16731_ ;
  assign \new_Sorter100|16832_  = \new_Sorter100|16732_  & \new_Sorter100|16733_ ;
  assign \new_Sorter100|16833_  = \new_Sorter100|16732_  | \new_Sorter100|16733_ ;
  assign \new_Sorter100|16834_  = \new_Sorter100|16734_  & \new_Sorter100|16735_ ;
  assign \new_Sorter100|16835_  = \new_Sorter100|16734_  | \new_Sorter100|16735_ ;
  assign \new_Sorter100|16836_  = \new_Sorter100|16736_  & \new_Sorter100|16737_ ;
  assign \new_Sorter100|16837_  = \new_Sorter100|16736_  | \new_Sorter100|16737_ ;
  assign \new_Sorter100|16838_  = \new_Sorter100|16738_  & \new_Sorter100|16739_ ;
  assign \new_Sorter100|16839_  = \new_Sorter100|16738_  | \new_Sorter100|16739_ ;
  assign \new_Sorter100|16840_  = \new_Sorter100|16740_  & \new_Sorter100|16741_ ;
  assign \new_Sorter100|16841_  = \new_Sorter100|16740_  | \new_Sorter100|16741_ ;
  assign \new_Sorter100|16842_  = \new_Sorter100|16742_  & \new_Sorter100|16743_ ;
  assign \new_Sorter100|16843_  = \new_Sorter100|16742_  | \new_Sorter100|16743_ ;
  assign \new_Sorter100|16844_  = \new_Sorter100|16744_  & \new_Sorter100|16745_ ;
  assign \new_Sorter100|16845_  = \new_Sorter100|16744_  | \new_Sorter100|16745_ ;
  assign \new_Sorter100|16846_  = \new_Sorter100|16746_  & \new_Sorter100|16747_ ;
  assign \new_Sorter100|16847_  = \new_Sorter100|16746_  | \new_Sorter100|16747_ ;
  assign \new_Sorter100|16848_  = \new_Sorter100|16748_  & \new_Sorter100|16749_ ;
  assign \new_Sorter100|16849_  = \new_Sorter100|16748_  | \new_Sorter100|16749_ ;
  assign \new_Sorter100|16850_  = \new_Sorter100|16750_  & \new_Sorter100|16751_ ;
  assign \new_Sorter100|16851_  = \new_Sorter100|16750_  | \new_Sorter100|16751_ ;
  assign \new_Sorter100|16852_  = \new_Sorter100|16752_  & \new_Sorter100|16753_ ;
  assign \new_Sorter100|16853_  = \new_Sorter100|16752_  | \new_Sorter100|16753_ ;
  assign \new_Sorter100|16854_  = \new_Sorter100|16754_  & \new_Sorter100|16755_ ;
  assign \new_Sorter100|16855_  = \new_Sorter100|16754_  | \new_Sorter100|16755_ ;
  assign \new_Sorter100|16856_  = \new_Sorter100|16756_  & \new_Sorter100|16757_ ;
  assign \new_Sorter100|16857_  = \new_Sorter100|16756_  | \new_Sorter100|16757_ ;
  assign \new_Sorter100|16858_  = \new_Sorter100|16758_  & \new_Sorter100|16759_ ;
  assign \new_Sorter100|16859_  = \new_Sorter100|16758_  | \new_Sorter100|16759_ ;
  assign \new_Sorter100|16860_  = \new_Sorter100|16760_  & \new_Sorter100|16761_ ;
  assign \new_Sorter100|16861_  = \new_Sorter100|16760_  | \new_Sorter100|16761_ ;
  assign \new_Sorter100|16862_  = \new_Sorter100|16762_  & \new_Sorter100|16763_ ;
  assign \new_Sorter100|16863_  = \new_Sorter100|16762_  | \new_Sorter100|16763_ ;
  assign \new_Sorter100|16864_  = \new_Sorter100|16764_  & \new_Sorter100|16765_ ;
  assign \new_Sorter100|16865_  = \new_Sorter100|16764_  | \new_Sorter100|16765_ ;
  assign \new_Sorter100|16866_  = \new_Sorter100|16766_  & \new_Sorter100|16767_ ;
  assign \new_Sorter100|16867_  = \new_Sorter100|16766_  | \new_Sorter100|16767_ ;
  assign \new_Sorter100|16868_  = \new_Sorter100|16768_  & \new_Sorter100|16769_ ;
  assign \new_Sorter100|16869_  = \new_Sorter100|16768_  | \new_Sorter100|16769_ ;
  assign \new_Sorter100|16870_  = \new_Sorter100|16770_  & \new_Sorter100|16771_ ;
  assign \new_Sorter100|16871_  = \new_Sorter100|16770_  | \new_Sorter100|16771_ ;
  assign \new_Sorter100|16872_  = \new_Sorter100|16772_  & \new_Sorter100|16773_ ;
  assign \new_Sorter100|16873_  = \new_Sorter100|16772_  | \new_Sorter100|16773_ ;
  assign \new_Sorter100|16874_  = \new_Sorter100|16774_  & \new_Sorter100|16775_ ;
  assign \new_Sorter100|16875_  = \new_Sorter100|16774_  | \new_Sorter100|16775_ ;
  assign \new_Sorter100|16876_  = \new_Sorter100|16776_  & \new_Sorter100|16777_ ;
  assign \new_Sorter100|16877_  = \new_Sorter100|16776_  | \new_Sorter100|16777_ ;
  assign \new_Sorter100|16878_  = \new_Sorter100|16778_  & \new_Sorter100|16779_ ;
  assign \new_Sorter100|16879_  = \new_Sorter100|16778_  | \new_Sorter100|16779_ ;
  assign \new_Sorter100|16880_  = \new_Sorter100|16780_  & \new_Sorter100|16781_ ;
  assign \new_Sorter100|16881_  = \new_Sorter100|16780_  | \new_Sorter100|16781_ ;
  assign \new_Sorter100|16882_  = \new_Sorter100|16782_  & \new_Sorter100|16783_ ;
  assign \new_Sorter100|16883_  = \new_Sorter100|16782_  | \new_Sorter100|16783_ ;
  assign \new_Sorter100|16884_  = \new_Sorter100|16784_  & \new_Sorter100|16785_ ;
  assign \new_Sorter100|16885_  = \new_Sorter100|16784_  | \new_Sorter100|16785_ ;
  assign \new_Sorter100|16886_  = \new_Sorter100|16786_  & \new_Sorter100|16787_ ;
  assign \new_Sorter100|16887_  = \new_Sorter100|16786_  | \new_Sorter100|16787_ ;
  assign \new_Sorter100|16888_  = \new_Sorter100|16788_  & \new_Sorter100|16789_ ;
  assign \new_Sorter100|16889_  = \new_Sorter100|16788_  | \new_Sorter100|16789_ ;
  assign \new_Sorter100|16890_  = \new_Sorter100|16790_  & \new_Sorter100|16791_ ;
  assign \new_Sorter100|16891_  = \new_Sorter100|16790_  | \new_Sorter100|16791_ ;
  assign \new_Sorter100|16892_  = \new_Sorter100|16792_  & \new_Sorter100|16793_ ;
  assign \new_Sorter100|16893_  = \new_Sorter100|16792_  | \new_Sorter100|16793_ ;
  assign \new_Sorter100|16894_  = \new_Sorter100|16794_  & \new_Sorter100|16795_ ;
  assign \new_Sorter100|16895_  = \new_Sorter100|16794_  | \new_Sorter100|16795_ ;
  assign \new_Sorter100|16896_  = \new_Sorter100|16796_  & \new_Sorter100|16797_ ;
  assign \new_Sorter100|16897_  = \new_Sorter100|16796_  | \new_Sorter100|16797_ ;
  assign \new_Sorter100|16898_  = \new_Sorter100|16798_  & \new_Sorter100|16799_ ;
  assign \new_Sorter100|16899_  = \new_Sorter100|16798_  | \new_Sorter100|16799_ ;
  assign \new_Sorter100|16900_  = \new_Sorter100|16800_ ;
  assign \new_Sorter100|16999_  = \new_Sorter100|16899_ ;
  assign \new_Sorter100|16901_  = \new_Sorter100|16801_  & \new_Sorter100|16802_ ;
  assign \new_Sorter100|16902_  = \new_Sorter100|16801_  | \new_Sorter100|16802_ ;
  assign \new_Sorter100|16903_  = \new_Sorter100|16803_  & \new_Sorter100|16804_ ;
  assign \new_Sorter100|16904_  = \new_Sorter100|16803_  | \new_Sorter100|16804_ ;
  assign \new_Sorter100|16905_  = \new_Sorter100|16805_  & \new_Sorter100|16806_ ;
  assign \new_Sorter100|16906_  = \new_Sorter100|16805_  | \new_Sorter100|16806_ ;
  assign \new_Sorter100|16907_  = \new_Sorter100|16807_  & \new_Sorter100|16808_ ;
  assign \new_Sorter100|16908_  = \new_Sorter100|16807_  | \new_Sorter100|16808_ ;
  assign \new_Sorter100|16909_  = \new_Sorter100|16809_  & \new_Sorter100|16810_ ;
  assign \new_Sorter100|16910_  = \new_Sorter100|16809_  | \new_Sorter100|16810_ ;
  assign \new_Sorter100|16911_  = \new_Sorter100|16811_  & \new_Sorter100|16812_ ;
  assign \new_Sorter100|16912_  = \new_Sorter100|16811_  | \new_Sorter100|16812_ ;
  assign \new_Sorter100|16913_  = \new_Sorter100|16813_  & \new_Sorter100|16814_ ;
  assign \new_Sorter100|16914_  = \new_Sorter100|16813_  | \new_Sorter100|16814_ ;
  assign \new_Sorter100|16915_  = \new_Sorter100|16815_  & \new_Sorter100|16816_ ;
  assign \new_Sorter100|16916_  = \new_Sorter100|16815_  | \new_Sorter100|16816_ ;
  assign \new_Sorter100|16917_  = \new_Sorter100|16817_  & \new_Sorter100|16818_ ;
  assign \new_Sorter100|16918_  = \new_Sorter100|16817_  | \new_Sorter100|16818_ ;
  assign \new_Sorter100|16919_  = \new_Sorter100|16819_  & \new_Sorter100|16820_ ;
  assign \new_Sorter100|16920_  = \new_Sorter100|16819_  | \new_Sorter100|16820_ ;
  assign \new_Sorter100|16921_  = \new_Sorter100|16821_  & \new_Sorter100|16822_ ;
  assign \new_Sorter100|16922_  = \new_Sorter100|16821_  | \new_Sorter100|16822_ ;
  assign \new_Sorter100|16923_  = \new_Sorter100|16823_  & \new_Sorter100|16824_ ;
  assign \new_Sorter100|16924_  = \new_Sorter100|16823_  | \new_Sorter100|16824_ ;
  assign \new_Sorter100|16925_  = \new_Sorter100|16825_  & \new_Sorter100|16826_ ;
  assign \new_Sorter100|16926_  = \new_Sorter100|16825_  | \new_Sorter100|16826_ ;
  assign \new_Sorter100|16927_  = \new_Sorter100|16827_  & \new_Sorter100|16828_ ;
  assign \new_Sorter100|16928_  = \new_Sorter100|16827_  | \new_Sorter100|16828_ ;
  assign \new_Sorter100|16929_  = \new_Sorter100|16829_  & \new_Sorter100|16830_ ;
  assign \new_Sorter100|16930_  = \new_Sorter100|16829_  | \new_Sorter100|16830_ ;
  assign \new_Sorter100|16931_  = \new_Sorter100|16831_  & \new_Sorter100|16832_ ;
  assign \new_Sorter100|16932_  = \new_Sorter100|16831_  | \new_Sorter100|16832_ ;
  assign \new_Sorter100|16933_  = \new_Sorter100|16833_  & \new_Sorter100|16834_ ;
  assign \new_Sorter100|16934_  = \new_Sorter100|16833_  | \new_Sorter100|16834_ ;
  assign \new_Sorter100|16935_  = \new_Sorter100|16835_  & \new_Sorter100|16836_ ;
  assign \new_Sorter100|16936_  = \new_Sorter100|16835_  | \new_Sorter100|16836_ ;
  assign \new_Sorter100|16937_  = \new_Sorter100|16837_  & \new_Sorter100|16838_ ;
  assign \new_Sorter100|16938_  = \new_Sorter100|16837_  | \new_Sorter100|16838_ ;
  assign \new_Sorter100|16939_  = \new_Sorter100|16839_  & \new_Sorter100|16840_ ;
  assign \new_Sorter100|16940_  = \new_Sorter100|16839_  | \new_Sorter100|16840_ ;
  assign \new_Sorter100|16941_  = \new_Sorter100|16841_  & \new_Sorter100|16842_ ;
  assign \new_Sorter100|16942_  = \new_Sorter100|16841_  | \new_Sorter100|16842_ ;
  assign \new_Sorter100|16943_  = \new_Sorter100|16843_  & \new_Sorter100|16844_ ;
  assign \new_Sorter100|16944_  = \new_Sorter100|16843_  | \new_Sorter100|16844_ ;
  assign \new_Sorter100|16945_  = \new_Sorter100|16845_  & \new_Sorter100|16846_ ;
  assign \new_Sorter100|16946_  = \new_Sorter100|16845_  | \new_Sorter100|16846_ ;
  assign \new_Sorter100|16947_  = \new_Sorter100|16847_  & \new_Sorter100|16848_ ;
  assign \new_Sorter100|16948_  = \new_Sorter100|16847_  | \new_Sorter100|16848_ ;
  assign \new_Sorter100|16949_  = \new_Sorter100|16849_  & \new_Sorter100|16850_ ;
  assign \new_Sorter100|16950_  = \new_Sorter100|16849_  | \new_Sorter100|16850_ ;
  assign \new_Sorter100|16951_  = \new_Sorter100|16851_  & \new_Sorter100|16852_ ;
  assign \new_Sorter100|16952_  = \new_Sorter100|16851_  | \new_Sorter100|16852_ ;
  assign \new_Sorter100|16953_  = \new_Sorter100|16853_  & \new_Sorter100|16854_ ;
  assign \new_Sorter100|16954_  = \new_Sorter100|16853_  | \new_Sorter100|16854_ ;
  assign \new_Sorter100|16955_  = \new_Sorter100|16855_  & \new_Sorter100|16856_ ;
  assign \new_Sorter100|16956_  = \new_Sorter100|16855_  | \new_Sorter100|16856_ ;
  assign \new_Sorter100|16957_  = \new_Sorter100|16857_  & \new_Sorter100|16858_ ;
  assign \new_Sorter100|16958_  = \new_Sorter100|16857_  | \new_Sorter100|16858_ ;
  assign \new_Sorter100|16959_  = \new_Sorter100|16859_  & \new_Sorter100|16860_ ;
  assign \new_Sorter100|16960_  = \new_Sorter100|16859_  | \new_Sorter100|16860_ ;
  assign \new_Sorter100|16961_  = \new_Sorter100|16861_  & \new_Sorter100|16862_ ;
  assign \new_Sorter100|16962_  = \new_Sorter100|16861_  | \new_Sorter100|16862_ ;
  assign \new_Sorter100|16963_  = \new_Sorter100|16863_  & \new_Sorter100|16864_ ;
  assign \new_Sorter100|16964_  = \new_Sorter100|16863_  | \new_Sorter100|16864_ ;
  assign \new_Sorter100|16965_  = \new_Sorter100|16865_  & \new_Sorter100|16866_ ;
  assign \new_Sorter100|16966_  = \new_Sorter100|16865_  | \new_Sorter100|16866_ ;
  assign \new_Sorter100|16967_  = \new_Sorter100|16867_  & \new_Sorter100|16868_ ;
  assign \new_Sorter100|16968_  = \new_Sorter100|16867_  | \new_Sorter100|16868_ ;
  assign \new_Sorter100|16969_  = \new_Sorter100|16869_  & \new_Sorter100|16870_ ;
  assign \new_Sorter100|16970_  = \new_Sorter100|16869_  | \new_Sorter100|16870_ ;
  assign \new_Sorter100|16971_  = \new_Sorter100|16871_  & \new_Sorter100|16872_ ;
  assign \new_Sorter100|16972_  = \new_Sorter100|16871_  | \new_Sorter100|16872_ ;
  assign \new_Sorter100|16973_  = \new_Sorter100|16873_  & \new_Sorter100|16874_ ;
  assign \new_Sorter100|16974_  = \new_Sorter100|16873_  | \new_Sorter100|16874_ ;
  assign \new_Sorter100|16975_  = \new_Sorter100|16875_  & \new_Sorter100|16876_ ;
  assign \new_Sorter100|16976_  = \new_Sorter100|16875_  | \new_Sorter100|16876_ ;
  assign \new_Sorter100|16977_  = \new_Sorter100|16877_  & \new_Sorter100|16878_ ;
  assign \new_Sorter100|16978_  = \new_Sorter100|16877_  | \new_Sorter100|16878_ ;
  assign \new_Sorter100|16979_  = \new_Sorter100|16879_  & \new_Sorter100|16880_ ;
  assign \new_Sorter100|16980_  = \new_Sorter100|16879_  | \new_Sorter100|16880_ ;
  assign \new_Sorter100|16981_  = \new_Sorter100|16881_  & \new_Sorter100|16882_ ;
  assign \new_Sorter100|16982_  = \new_Sorter100|16881_  | \new_Sorter100|16882_ ;
  assign \new_Sorter100|16983_  = \new_Sorter100|16883_  & \new_Sorter100|16884_ ;
  assign \new_Sorter100|16984_  = \new_Sorter100|16883_  | \new_Sorter100|16884_ ;
  assign \new_Sorter100|16985_  = \new_Sorter100|16885_  & \new_Sorter100|16886_ ;
  assign \new_Sorter100|16986_  = \new_Sorter100|16885_  | \new_Sorter100|16886_ ;
  assign \new_Sorter100|16987_  = \new_Sorter100|16887_  & \new_Sorter100|16888_ ;
  assign \new_Sorter100|16988_  = \new_Sorter100|16887_  | \new_Sorter100|16888_ ;
  assign \new_Sorter100|16989_  = \new_Sorter100|16889_  & \new_Sorter100|16890_ ;
  assign \new_Sorter100|16990_  = \new_Sorter100|16889_  | \new_Sorter100|16890_ ;
  assign \new_Sorter100|16991_  = \new_Sorter100|16891_  & \new_Sorter100|16892_ ;
  assign \new_Sorter100|16992_  = \new_Sorter100|16891_  | \new_Sorter100|16892_ ;
  assign \new_Sorter100|16993_  = \new_Sorter100|16893_  & \new_Sorter100|16894_ ;
  assign \new_Sorter100|16994_  = \new_Sorter100|16893_  | \new_Sorter100|16894_ ;
  assign \new_Sorter100|16995_  = \new_Sorter100|16895_  & \new_Sorter100|16896_ ;
  assign \new_Sorter100|16996_  = \new_Sorter100|16895_  | \new_Sorter100|16896_ ;
  assign \new_Sorter100|16997_  = \new_Sorter100|16897_  & \new_Sorter100|16898_ ;
  assign \new_Sorter100|16998_  = \new_Sorter100|16897_  | \new_Sorter100|16898_ ;
  assign \new_Sorter100|17000_  = \new_Sorter100|16900_  & \new_Sorter100|16901_ ;
  assign \new_Sorter100|17001_  = \new_Sorter100|16900_  | \new_Sorter100|16901_ ;
  assign \new_Sorter100|17002_  = \new_Sorter100|16902_  & \new_Sorter100|16903_ ;
  assign \new_Sorter100|17003_  = \new_Sorter100|16902_  | \new_Sorter100|16903_ ;
  assign \new_Sorter100|17004_  = \new_Sorter100|16904_  & \new_Sorter100|16905_ ;
  assign \new_Sorter100|17005_  = \new_Sorter100|16904_  | \new_Sorter100|16905_ ;
  assign \new_Sorter100|17006_  = \new_Sorter100|16906_  & \new_Sorter100|16907_ ;
  assign \new_Sorter100|17007_  = \new_Sorter100|16906_  | \new_Sorter100|16907_ ;
  assign \new_Sorter100|17008_  = \new_Sorter100|16908_  & \new_Sorter100|16909_ ;
  assign \new_Sorter100|17009_  = \new_Sorter100|16908_  | \new_Sorter100|16909_ ;
  assign \new_Sorter100|17010_  = \new_Sorter100|16910_  & \new_Sorter100|16911_ ;
  assign \new_Sorter100|17011_  = \new_Sorter100|16910_  | \new_Sorter100|16911_ ;
  assign \new_Sorter100|17012_  = \new_Sorter100|16912_  & \new_Sorter100|16913_ ;
  assign \new_Sorter100|17013_  = \new_Sorter100|16912_  | \new_Sorter100|16913_ ;
  assign \new_Sorter100|17014_  = \new_Sorter100|16914_  & \new_Sorter100|16915_ ;
  assign \new_Sorter100|17015_  = \new_Sorter100|16914_  | \new_Sorter100|16915_ ;
  assign \new_Sorter100|17016_  = \new_Sorter100|16916_  & \new_Sorter100|16917_ ;
  assign \new_Sorter100|17017_  = \new_Sorter100|16916_  | \new_Sorter100|16917_ ;
  assign \new_Sorter100|17018_  = \new_Sorter100|16918_  & \new_Sorter100|16919_ ;
  assign \new_Sorter100|17019_  = \new_Sorter100|16918_  | \new_Sorter100|16919_ ;
  assign \new_Sorter100|17020_  = \new_Sorter100|16920_  & \new_Sorter100|16921_ ;
  assign \new_Sorter100|17021_  = \new_Sorter100|16920_  | \new_Sorter100|16921_ ;
  assign \new_Sorter100|17022_  = \new_Sorter100|16922_  & \new_Sorter100|16923_ ;
  assign \new_Sorter100|17023_  = \new_Sorter100|16922_  | \new_Sorter100|16923_ ;
  assign \new_Sorter100|17024_  = \new_Sorter100|16924_  & \new_Sorter100|16925_ ;
  assign \new_Sorter100|17025_  = \new_Sorter100|16924_  | \new_Sorter100|16925_ ;
  assign \new_Sorter100|17026_  = \new_Sorter100|16926_  & \new_Sorter100|16927_ ;
  assign \new_Sorter100|17027_  = \new_Sorter100|16926_  | \new_Sorter100|16927_ ;
  assign \new_Sorter100|17028_  = \new_Sorter100|16928_  & \new_Sorter100|16929_ ;
  assign \new_Sorter100|17029_  = \new_Sorter100|16928_  | \new_Sorter100|16929_ ;
  assign \new_Sorter100|17030_  = \new_Sorter100|16930_  & \new_Sorter100|16931_ ;
  assign \new_Sorter100|17031_  = \new_Sorter100|16930_  | \new_Sorter100|16931_ ;
  assign \new_Sorter100|17032_  = \new_Sorter100|16932_  & \new_Sorter100|16933_ ;
  assign \new_Sorter100|17033_  = \new_Sorter100|16932_  | \new_Sorter100|16933_ ;
  assign \new_Sorter100|17034_  = \new_Sorter100|16934_  & \new_Sorter100|16935_ ;
  assign \new_Sorter100|17035_  = \new_Sorter100|16934_  | \new_Sorter100|16935_ ;
  assign \new_Sorter100|17036_  = \new_Sorter100|16936_  & \new_Sorter100|16937_ ;
  assign \new_Sorter100|17037_  = \new_Sorter100|16936_  | \new_Sorter100|16937_ ;
  assign \new_Sorter100|17038_  = \new_Sorter100|16938_  & \new_Sorter100|16939_ ;
  assign \new_Sorter100|17039_  = \new_Sorter100|16938_  | \new_Sorter100|16939_ ;
  assign \new_Sorter100|17040_  = \new_Sorter100|16940_  & \new_Sorter100|16941_ ;
  assign \new_Sorter100|17041_  = \new_Sorter100|16940_  | \new_Sorter100|16941_ ;
  assign \new_Sorter100|17042_  = \new_Sorter100|16942_  & \new_Sorter100|16943_ ;
  assign \new_Sorter100|17043_  = \new_Sorter100|16942_  | \new_Sorter100|16943_ ;
  assign \new_Sorter100|17044_  = \new_Sorter100|16944_  & \new_Sorter100|16945_ ;
  assign \new_Sorter100|17045_  = \new_Sorter100|16944_  | \new_Sorter100|16945_ ;
  assign \new_Sorter100|17046_  = \new_Sorter100|16946_  & \new_Sorter100|16947_ ;
  assign \new_Sorter100|17047_  = \new_Sorter100|16946_  | \new_Sorter100|16947_ ;
  assign \new_Sorter100|17048_  = \new_Sorter100|16948_  & \new_Sorter100|16949_ ;
  assign \new_Sorter100|17049_  = \new_Sorter100|16948_  | \new_Sorter100|16949_ ;
  assign \new_Sorter100|17050_  = \new_Sorter100|16950_  & \new_Sorter100|16951_ ;
  assign \new_Sorter100|17051_  = \new_Sorter100|16950_  | \new_Sorter100|16951_ ;
  assign \new_Sorter100|17052_  = \new_Sorter100|16952_  & \new_Sorter100|16953_ ;
  assign \new_Sorter100|17053_  = \new_Sorter100|16952_  | \new_Sorter100|16953_ ;
  assign \new_Sorter100|17054_  = \new_Sorter100|16954_  & \new_Sorter100|16955_ ;
  assign \new_Sorter100|17055_  = \new_Sorter100|16954_  | \new_Sorter100|16955_ ;
  assign \new_Sorter100|17056_  = \new_Sorter100|16956_  & \new_Sorter100|16957_ ;
  assign \new_Sorter100|17057_  = \new_Sorter100|16956_  | \new_Sorter100|16957_ ;
  assign \new_Sorter100|17058_  = \new_Sorter100|16958_  & \new_Sorter100|16959_ ;
  assign \new_Sorter100|17059_  = \new_Sorter100|16958_  | \new_Sorter100|16959_ ;
  assign \new_Sorter100|17060_  = \new_Sorter100|16960_  & \new_Sorter100|16961_ ;
  assign \new_Sorter100|17061_  = \new_Sorter100|16960_  | \new_Sorter100|16961_ ;
  assign \new_Sorter100|17062_  = \new_Sorter100|16962_  & \new_Sorter100|16963_ ;
  assign \new_Sorter100|17063_  = \new_Sorter100|16962_  | \new_Sorter100|16963_ ;
  assign \new_Sorter100|17064_  = \new_Sorter100|16964_  & \new_Sorter100|16965_ ;
  assign \new_Sorter100|17065_  = \new_Sorter100|16964_  | \new_Sorter100|16965_ ;
  assign \new_Sorter100|17066_  = \new_Sorter100|16966_  & \new_Sorter100|16967_ ;
  assign \new_Sorter100|17067_  = \new_Sorter100|16966_  | \new_Sorter100|16967_ ;
  assign \new_Sorter100|17068_  = \new_Sorter100|16968_  & \new_Sorter100|16969_ ;
  assign \new_Sorter100|17069_  = \new_Sorter100|16968_  | \new_Sorter100|16969_ ;
  assign \new_Sorter100|17070_  = \new_Sorter100|16970_  & \new_Sorter100|16971_ ;
  assign \new_Sorter100|17071_  = \new_Sorter100|16970_  | \new_Sorter100|16971_ ;
  assign \new_Sorter100|17072_  = \new_Sorter100|16972_  & \new_Sorter100|16973_ ;
  assign \new_Sorter100|17073_  = \new_Sorter100|16972_  | \new_Sorter100|16973_ ;
  assign \new_Sorter100|17074_  = \new_Sorter100|16974_  & \new_Sorter100|16975_ ;
  assign \new_Sorter100|17075_  = \new_Sorter100|16974_  | \new_Sorter100|16975_ ;
  assign \new_Sorter100|17076_  = \new_Sorter100|16976_  & \new_Sorter100|16977_ ;
  assign \new_Sorter100|17077_  = \new_Sorter100|16976_  | \new_Sorter100|16977_ ;
  assign \new_Sorter100|17078_  = \new_Sorter100|16978_  & \new_Sorter100|16979_ ;
  assign \new_Sorter100|17079_  = \new_Sorter100|16978_  | \new_Sorter100|16979_ ;
  assign \new_Sorter100|17080_  = \new_Sorter100|16980_  & \new_Sorter100|16981_ ;
  assign \new_Sorter100|17081_  = \new_Sorter100|16980_  | \new_Sorter100|16981_ ;
  assign \new_Sorter100|17082_  = \new_Sorter100|16982_  & \new_Sorter100|16983_ ;
  assign \new_Sorter100|17083_  = \new_Sorter100|16982_  | \new_Sorter100|16983_ ;
  assign \new_Sorter100|17084_  = \new_Sorter100|16984_  & \new_Sorter100|16985_ ;
  assign \new_Sorter100|17085_  = \new_Sorter100|16984_  | \new_Sorter100|16985_ ;
  assign \new_Sorter100|17086_  = \new_Sorter100|16986_  & \new_Sorter100|16987_ ;
  assign \new_Sorter100|17087_  = \new_Sorter100|16986_  | \new_Sorter100|16987_ ;
  assign \new_Sorter100|17088_  = \new_Sorter100|16988_  & \new_Sorter100|16989_ ;
  assign \new_Sorter100|17089_  = \new_Sorter100|16988_  | \new_Sorter100|16989_ ;
  assign \new_Sorter100|17090_  = \new_Sorter100|16990_  & \new_Sorter100|16991_ ;
  assign \new_Sorter100|17091_  = \new_Sorter100|16990_  | \new_Sorter100|16991_ ;
  assign \new_Sorter100|17092_  = \new_Sorter100|16992_  & \new_Sorter100|16993_ ;
  assign \new_Sorter100|17093_  = \new_Sorter100|16992_  | \new_Sorter100|16993_ ;
  assign \new_Sorter100|17094_  = \new_Sorter100|16994_  & \new_Sorter100|16995_ ;
  assign \new_Sorter100|17095_  = \new_Sorter100|16994_  | \new_Sorter100|16995_ ;
  assign \new_Sorter100|17096_  = \new_Sorter100|16996_  & \new_Sorter100|16997_ ;
  assign \new_Sorter100|17097_  = \new_Sorter100|16996_  | \new_Sorter100|16997_ ;
  assign \new_Sorter100|17098_  = \new_Sorter100|16998_  & \new_Sorter100|16999_ ;
  assign \new_Sorter100|17099_  = \new_Sorter100|16998_  | \new_Sorter100|16999_ ;
  assign \new_Sorter100|17100_  = \new_Sorter100|17000_ ;
  assign \new_Sorter100|17199_  = \new_Sorter100|17099_ ;
  assign \new_Sorter100|17101_  = \new_Sorter100|17001_  & \new_Sorter100|17002_ ;
  assign \new_Sorter100|17102_  = \new_Sorter100|17001_  | \new_Sorter100|17002_ ;
  assign \new_Sorter100|17103_  = \new_Sorter100|17003_  & \new_Sorter100|17004_ ;
  assign \new_Sorter100|17104_  = \new_Sorter100|17003_  | \new_Sorter100|17004_ ;
  assign \new_Sorter100|17105_  = \new_Sorter100|17005_  & \new_Sorter100|17006_ ;
  assign \new_Sorter100|17106_  = \new_Sorter100|17005_  | \new_Sorter100|17006_ ;
  assign \new_Sorter100|17107_  = \new_Sorter100|17007_  & \new_Sorter100|17008_ ;
  assign \new_Sorter100|17108_  = \new_Sorter100|17007_  | \new_Sorter100|17008_ ;
  assign \new_Sorter100|17109_  = \new_Sorter100|17009_  & \new_Sorter100|17010_ ;
  assign \new_Sorter100|17110_  = \new_Sorter100|17009_  | \new_Sorter100|17010_ ;
  assign \new_Sorter100|17111_  = \new_Sorter100|17011_  & \new_Sorter100|17012_ ;
  assign \new_Sorter100|17112_  = \new_Sorter100|17011_  | \new_Sorter100|17012_ ;
  assign \new_Sorter100|17113_  = \new_Sorter100|17013_  & \new_Sorter100|17014_ ;
  assign \new_Sorter100|17114_  = \new_Sorter100|17013_  | \new_Sorter100|17014_ ;
  assign \new_Sorter100|17115_  = \new_Sorter100|17015_  & \new_Sorter100|17016_ ;
  assign \new_Sorter100|17116_  = \new_Sorter100|17015_  | \new_Sorter100|17016_ ;
  assign \new_Sorter100|17117_  = \new_Sorter100|17017_  & \new_Sorter100|17018_ ;
  assign \new_Sorter100|17118_  = \new_Sorter100|17017_  | \new_Sorter100|17018_ ;
  assign \new_Sorter100|17119_  = \new_Sorter100|17019_  & \new_Sorter100|17020_ ;
  assign \new_Sorter100|17120_  = \new_Sorter100|17019_  | \new_Sorter100|17020_ ;
  assign \new_Sorter100|17121_  = \new_Sorter100|17021_  & \new_Sorter100|17022_ ;
  assign \new_Sorter100|17122_  = \new_Sorter100|17021_  | \new_Sorter100|17022_ ;
  assign \new_Sorter100|17123_  = \new_Sorter100|17023_  & \new_Sorter100|17024_ ;
  assign \new_Sorter100|17124_  = \new_Sorter100|17023_  | \new_Sorter100|17024_ ;
  assign \new_Sorter100|17125_  = \new_Sorter100|17025_  & \new_Sorter100|17026_ ;
  assign \new_Sorter100|17126_  = \new_Sorter100|17025_  | \new_Sorter100|17026_ ;
  assign \new_Sorter100|17127_  = \new_Sorter100|17027_  & \new_Sorter100|17028_ ;
  assign \new_Sorter100|17128_  = \new_Sorter100|17027_  | \new_Sorter100|17028_ ;
  assign \new_Sorter100|17129_  = \new_Sorter100|17029_  & \new_Sorter100|17030_ ;
  assign \new_Sorter100|17130_  = \new_Sorter100|17029_  | \new_Sorter100|17030_ ;
  assign \new_Sorter100|17131_  = \new_Sorter100|17031_  & \new_Sorter100|17032_ ;
  assign \new_Sorter100|17132_  = \new_Sorter100|17031_  | \new_Sorter100|17032_ ;
  assign \new_Sorter100|17133_  = \new_Sorter100|17033_  & \new_Sorter100|17034_ ;
  assign \new_Sorter100|17134_  = \new_Sorter100|17033_  | \new_Sorter100|17034_ ;
  assign \new_Sorter100|17135_  = \new_Sorter100|17035_  & \new_Sorter100|17036_ ;
  assign \new_Sorter100|17136_  = \new_Sorter100|17035_  | \new_Sorter100|17036_ ;
  assign \new_Sorter100|17137_  = \new_Sorter100|17037_  & \new_Sorter100|17038_ ;
  assign \new_Sorter100|17138_  = \new_Sorter100|17037_  | \new_Sorter100|17038_ ;
  assign \new_Sorter100|17139_  = \new_Sorter100|17039_  & \new_Sorter100|17040_ ;
  assign \new_Sorter100|17140_  = \new_Sorter100|17039_  | \new_Sorter100|17040_ ;
  assign \new_Sorter100|17141_  = \new_Sorter100|17041_  & \new_Sorter100|17042_ ;
  assign \new_Sorter100|17142_  = \new_Sorter100|17041_  | \new_Sorter100|17042_ ;
  assign \new_Sorter100|17143_  = \new_Sorter100|17043_  & \new_Sorter100|17044_ ;
  assign \new_Sorter100|17144_  = \new_Sorter100|17043_  | \new_Sorter100|17044_ ;
  assign \new_Sorter100|17145_  = \new_Sorter100|17045_  & \new_Sorter100|17046_ ;
  assign \new_Sorter100|17146_  = \new_Sorter100|17045_  | \new_Sorter100|17046_ ;
  assign \new_Sorter100|17147_  = \new_Sorter100|17047_  & \new_Sorter100|17048_ ;
  assign \new_Sorter100|17148_  = \new_Sorter100|17047_  | \new_Sorter100|17048_ ;
  assign \new_Sorter100|17149_  = \new_Sorter100|17049_  & \new_Sorter100|17050_ ;
  assign \new_Sorter100|17150_  = \new_Sorter100|17049_  | \new_Sorter100|17050_ ;
  assign \new_Sorter100|17151_  = \new_Sorter100|17051_  & \new_Sorter100|17052_ ;
  assign \new_Sorter100|17152_  = \new_Sorter100|17051_  | \new_Sorter100|17052_ ;
  assign \new_Sorter100|17153_  = \new_Sorter100|17053_  & \new_Sorter100|17054_ ;
  assign \new_Sorter100|17154_  = \new_Sorter100|17053_  | \new_Sorter100|17054_ ;
  assign \new_Sorter100|17155_  = \new_Sorter100|17055_  & \new_Sorter100|17056_ ;
  assign \new_Sorter100|17156_  = \new_Sorter100|17055_  | \new_Sorter100|17056_ ;
  assign \new_Sorter100|17157_  = \new_Sorter100|17057_  & \new_Sorter100|17058_ ;
  assign \new_Sorter100|17158_  = \new_Sorter100|17057_  | \new_Sorter100|17058_ ;
  assign \new_Sorter100|17159_  = \new_Sorter100|17059_  & \new_Sorter100|17060_ ;
  assign \new_Sorter100|17160_  = \new_Sorter100|17059_  | \new_Sorter100|17060_ ;
  assign \new_Sorter100|17161_  = \new_Sorter100|17061_  & \new_Sorter100|17062_ ;
  assign \new_Sorter100|17162_  = \new_Sorter100|17061_  | \new_Sorter100|17062_ ;
  assign \new_Sorter100|17163_  = \new_Sorter100|17063_  & \new_Sorter100|17064_ ;
  assign \new_Sorter100|17164_  = \new_Sorter100|17063_  | \new_Sorter100|17064_ ;
  assign \new_Sorter100|17165_  = \new_Sorter100|17065_  & \new_Sorter100|17066_ ;
  assign \new_Sorter100|17166_  = \new_Sorter100|17065_  | \new_Sorter100|17066_ ;
  assign \new_Sorter100|17167_  = \new_Sorter100|17067_  & \new_Sorter100|17068_ ;
  assign \new_Sorter100|17168_  = \new_Sorter100|17067_  | \new_Sorter100|17068_ ;
  assign \new_Sorter100|17169_  = \new_Sorter100|17069_  & \new_Sorter100|17070_ ;
  assign \new_Sorter100|17170_  = \new_Sorter100|17069_  | \new_Sorter100|17070_ ;
  assign \new_Sorter100|17171_  = \new_Sorter100|17071_  & \new_Sorter100|17072_ ;
  assign \new_Sorter100|17172_  = \new_Sorter100|17071_  | \new_Sorter100|17072_ ;
  assign \new_Sorter100|17173_  = \new_Sorter100|17073_  & \new_Sorter100|17074_ ;
  assign \new_Sorter100|17174_  = \new_Sorter100|17073_  | \new_Sorter100|17074_ ;
  assign \new_Sorter100|17175_  = \new_Sorter100|17075_  & \new_Sorter100|17076_ ;
  assign \new_Sorter100|17176_  = \new_Sorter100|17075_  | \new_Sorter100|17076_ ;
  assign \new_Sorter100|17177_  = \new_Sorter100|17077_  & \new_Sorter100|17078_ ;
  assign \new_Sorter100|17178_  = \new_Sorter100|17077_  | \new_Sorter100|17078_ ;
  assign \new_Sorter100|17179_  = \new_Sorter100|17079_  & \new_Sorter100|17080_ ;
  assign \new_Sorter100|17180_  = \new_Sorter100|17079_  | \new_Sorter100|17080_ ;
  assign \new_Sorter100|17181_  = \new_Sorter100|17081_  & \new_Sorter100|17082_ ;
  assign \new_Sorter100|17182_  = \new_Sorter100|17081_  | \new_Sorter100|17082_ ;
  assign \new_Sorter100|17183_  = \new_Sorter100|17083_  & \new_Sorter100|17084_ ;
  assign \new_Sorter100|17184_  = \new_Sorter100|17083_  | \new_Sorter100|17084_ ;
  assign \new_Sorter100|17185_  = \new_Sorter100|17085_  & \new_Sorter100|17086_ ;
  assign \new_Sorter100|17186_  = \new_Sorter100|17085_  | \new_Sorter100|17086_ ;
  assign \new_Sorter100|17187_  = \new_Sorter100|17087_  & \new_Sorter100|17088_ ;
  assign \new_Sorter100|17188_  = \new_Sorter100|17087_  | \new_Sorter100|17088_ ;
  assign \new_Sorter100|17189_  = \new_Sorter100|17089_  & \new_Sorter100|17090_ ;
  assign \new_Sorter100|17190_  = \new_Sorter100|17089_  | \new_Sorter100|17090_ ;
  assign \new_Sorter100|17191_  = \new_Sorter100|17091_  & \new_Sorter100|17092_ ;
  assign \new_Sorter100|17192_  = \new_Sorter100|17091_  | \new_Sorter100|17092_ ;
  assign \new_Sorter100|17193_  = \new_Sorter100|17093_  & \new_Sorter100|17094_ ;
  assign \new_Sorter100|17194_  = \new_Sorter100|17093_  | \new_Sorter100|17094_ ;
  assign \new_Sorter100|17195_  = \new_Sorter100|17095_  & \new_Sorter100|17096_ ;
  assign \new_Sorter100|17196_  = \new_Sorter100|17095_  | \new_Sorter100|17096_ ;
  assign \new_Sorter100|17197_  = \new_Sorter100|17097_  & \new_Sorter100|17098_ ;
  assign \new_Sorter100|17198_  = \new_Sorter100|17097_  | \new_Sorter100|17098_ ;
  assign \new_Sorter100|17200_  = \new_Sorter100|17100_  & \new_Sorter100|17101_ ;
  assign \new_Sorter100|17201_  = \new_Sorter100|17100_  | \new_Sorter100|17101_ ;
  assign \new_Sorter100|17202_  = \new_Sorter100|17102_  & \new_Sorter100|17103_ ;
  assign \new_Sorter100|17203_  = \new_Sorter100|17102_  | \new_Sorter100|17103_ ;
  assign \new_Sorter100|17204_  = \new_Sorter100|17104_  & \new_Sorter100|17105_ ;
  assign \new_Sorter100|17205_  = \new_Sorter100|17104_  | \new_Sorter100|17105_ ;
  assign \new_Sorter100|17206_  = \new_Sorter100|17106_  & \new_Sorter100|17107_ ;
  assign \new_Sorter100|17207_  = \new_Sorter100|17106_  | \new_Sorter100|17107_ ;
  assign \new_Sorter100|17208_  = \new_Sorter100|17108_  & \new_Sorter100|17109_ ;
  assign \new_Sorter100|17209_  = \new_Sorter100|17108_  | \new_Sorter100|17109_ ;
  assign \new_Sorter100|17210_  = \new_Sorter100|17110_  & \new_Sorter100|17111_ ;
  assign \new_Sorter100|17211_  = \new_Sorter100|17110_  | \new_Sorter100|17111_ ;
  assign \new_Sorter100|17212_  = \new_Sorter100|17112_  & \new_Sorter100|17113_ ;
  assign \new_Sorter100|17213_  = \new_Sorter100|17112_  | \new_Sorter100|17113_ ;
  assign \new_Sorter100|17214_  = \new_Sorter100|17114_  & \new_Sorter100|17115_ ;
  assign \new_Sorter100|17215_  = \new_Sorter100|17114_  | \new_Sorter100|17115_ ;
  assign \new_Sorter100|17216_  = \new_Sorter100|17116_  & \new_Sorter100|17117_ ;
  assign \new_Sorter100|17217_  = \new_Sorter100|17116_  | \new_Sorter100|17117_ ;
  assign \new_Sorter100|17218_  = \new_Sorter100|17118_  & \new_Sorter100|17119_ ;
  assign \new_Sorter100|17219_  = \new_Sorter100|17118_  | \new_Sorter100|17119_ ;
  assign \new_Sorter100|17220_  = \new_Sorter100|17120_  & \new_Sorter100|17121_ ;
  assign \new_Sorter100|17221_  = \new_Sorter100|17120_  | \new_Sorter100|17121_ ;
  assign \new_Sorter100|17222_  = \new_Sorter100|17122_  & \new_Sorter100|17123_ ;
  assign \new_Sorter100|17223_  = \new_Sorter100|17122_  | \new_Sorter100|17123_ ;
  assign \new_Sorter100|17224_  = \new_Sorter100|17124_  & \new_Sorter100|17125_ ;
  assign \new_Sorter100|17225_  = \new_Sorter100|17124_  | \new_Sorter100|17125_ ;
  assign \new_Sorter100|17226_  = \new_Sorter100|17126_  & \new_Sorter100|17127_ ;
  assign \new_Sorter100|17227_  = \new_Sorter100|17126_  | \new_Sorter100|17127_ ;
  assign \new_Sorter100|17228_  = \new_Sorter100|17128_  & \new_Sorter100|17129_ ;
  assign \new_Sorter100|17229_  = \new_Sorter100|17128_  | \new_Sorter100|17129_ ;
  assign \new_Sorter100|17230_  = \new_Sorter100|17130_  & \new_Sorter100|17131_ ;
  assign \new_Sorter100|17231_  = \new_Sorter100|17130_  | \new_Sorter100|17131_ ;
  assign \new_Sorter100|17232_  = \new_Sorter100|17132_  & \new_Sorter100|17133_ ;
  assign \new_Sorter100|17233_  = \new_Sorter100|17132_  | \new_Sorter100|17133_ ;
  assign \new_Sorter100|17234_  = \new_Sorter100|17134_  & \new_Sorter100|17135_ ;
  assign \new_Sorter100|17235_  = \new_Sorter100|17134_  | \new_Sorter100|17135_ ;
  assign \new_Sorter100|17236_  = \new_Sorter100|17136_  & \new_Sorter100|17137_ ;
  assign \new_Sorter100|17237_  = \new_Sorter100|17136_  | \new_Sorter100|17137_ ;
  assign \new_Sorter100|17238_  = \new_Sorter100|17138_  & \new_Sorter100|17139_ ;
  assign \new_Sorter100|17239_  = \new_Sorter100|17138_  | \new_Sorter100|17139_ ;
  assign \new_Sorter100|17240_  = \new_Sorter100|17140_  & \new_Sorter100|17141_ ;
  assign \new_Sorter100|17241_  = \new_Sorter100|17140_  | \new_Sorter100|17141_ ;
  assign \new_Sorter100|17242_  = \new_Sorter100|17142_  & \new_Sorter100|17143_ ;
  assign \new_Sorter100|17243_  = \new_Sorter100|17142_  | \new_Sorter100|17143_ ;
  assign \new_Sorter100|17244_  = \new_Sorter100|17144_  & \new_Sorter100|17145_ ;
  assign \new_Sorter100|17245_  = \new_Sorter100|17144_  | \new_Sorter100|17145_ ;
  assign \new_Sorter100|17246_  = \new_Sorter100|17146_  & \new_Sorter100|17147_ ;
  assign \new_Sorter100|17247_  = \new_Sorter100|17146_  | \new_Sorter100|17147_ ;
  assign \new_Sorter100|17248_  = \new_Sorter100|17148_  & \new_Sorter100|17149_ ;
  assign \new_Sorter100|17249_  = \new_Sorter100|17148_  | \new_Sorter100|17149_ ;
  assign \new_Sorter100|17250_  = \new_Sorter100|17150_  & \new_Sorter100|17151_ ;
  assign \new_Sorter100|17251_  = \new_Sorter100|17150_  | \new_Sorter100|17151_ ;
  assign \new_Sorter100|17252_  = \new_Sorter100|17152_  & \new_Sorter100|17153_ ;
  assign \new_Sorter100|17253_  = \new_Sorter100|17152_  | \new_Sorter100|17153_ ;
  assign \new_Sorter100|17254_  = \new_Sorter100|17154_  & \new_Sorter100|17155_ ;
  assign \new_Sorter100|17255_  = \new_Sorter100|17154_  | \new_Sorter100|17155_ ;
  assign \new_Sorter100|17256_  = \new_Sorter100|17156_  & \new_Sorter100|17157_ ;
  assign \new_Sorter100|17257_  = \new_Sorter100|17156_  | \new_Sorter100|17157_ ;
  assign \new_Sorter100|17258_  = \new_Sorter100|17158_  & \new_Sorter100|17159_ ;
  assign \new_Sorter100|17259_  = \new_Sorter100|17158_  | \new_Sorter100|17159_ ;
  assign \new_Sorter100|17260_  = \new_Sorter100|17160_  & \new_Sorter100|17161_ ;
  assign \new_Sorter100|17261_  = \new_Sorter100|17160_  | \new_Sorter100|17161_ ;
  assign \new_Sorter100|17262_  = \new_Sorter100|17162_  & \new_Sorter100|17163_ ;
  assign \new_Sorter100|17263_  = \new_Sorter100|17162_  | \new_Sorter100|17163_ ;
  assign \new_Sorter100|17264_  = \new_Sorter100|17164_  & \new_Sorter100|17165_ ;
  assign \new_Sorter100|17265_  = \new_Sorter100|17164_  | \new_Sorter100|17165_ ;
  assign \new_Sorter100|17266_  = \new_Sorter100|17166_  & \new_Sorter100|17167_ ;
  assign \new_Sorter100|17267_  = \new_Sorter100|17166_  | \new_Sorter100|17167_ ;
  assign \new_Sorter100|17268_  = \new_Sorter100|17168_  & \new_Sorter100|17169_ ;
  assign \new_Sorter100|17269_  = \new_Sorter100|17168_  | \new_Sorter100|17169_ ;
  assign \new_Sorter100|17270_  = \new_Sorter100|17170_  & \new_Sorter100|17171_ ;
  assign \new_Sorter100|17271_  = \new_Sorter100|17170_  | \new_Sorter100|17171_ ;
  assign \new_Sorter100|17272_  = \new_Sorter100|17172_  & \new_Sorter100|17173_ ;
  assign \new_Sorter100|17273_  = \new_Sorter100|17172_  | \new_Sorter100|17173_ ;
  assign \new_Sorter100|17274_  = \new_Sorter100|17174_  & \new_Sorter100|17175_ ;
  assign \new_Sorter100|17275_  = \new_Sorter100|17174_  | \new_Sorter100|17175_ ;
  assign \new_Sorter100|17276_  = \new_Sorter100|17176_  & \new_Sorter100|17177_ ;
  assign \new_Sorter100|17277_  = \new_Sorter100|17176_  | \new_Sorter100|17177_ ;
  assign \new_Sorter100|17278_  = \new_Sorter100|17178_  & \new_Sorter100|17179_ ;
  assign \new_Sorter100|17279_  = \new_Sorter100|17178_  | \new_Sorter100|17179_ ;
  assign \new_Sorter100|17280_  = \new_Sorter100|17180_  & \new_Sorter100|17181_ ;
  assign \new_Sorter100|17281_  = \new_Sorter100|17180_  | \new_Sorter100|17181_ ;
  assign \new_Sorter100|17282_  = \new_Sorter100|17182_  & \new_Sorter100|17183_ ;
  assign \new_Sorter100|17283_  = \new_Sorter100|17182_  | \new_Sorter100|17183_ ;
  assign \new_Sorter100|17284_  = \new_Sorter100|17184_  & \new_Sorter100|17185_ ;
  assign \new_Sorter100|17285_  = \new_Sorter100|17184_  | \new_Sorter100|17185_ ;
  assign \new_Sorter100|17286_  = \new_Sorter100|17186_  & \new_Sorter100|17187_ ;
  assign \new_Sorter100|17287_  = \new_Sorter100|17186_  | \new_Sorter100|17187_ ;
  assign \new_Sorter100|17288_  = \new_Sorter100|17188_  & \new_Sorter100|17189_ ;
  assign \new_Sorter100|17289_  = \new_Sorter100|17188_  | \new_Sorter100|17189_ ;
  assign \new_Sorter100|17290_  = \new_Sorter100|17190_  & \new_Sorter100|17191_ ;
  assign \new_Sorter100|17291_  = \new_Sorter100|17190_  | \new_Sorter100|17191_ ;
  assign \new_Sorter100|17292_  = \new_Sorter100|17192_  & \new_Sorter100|17193_ ;
  assign \new_Sorter100|17293_  = \new_Sorter100|17192_  | \new_Sorter100|17193_ ;
  assign \new_Sorter100|17294_  = \new_Sorter100|17194_  & \new_Sorter100|17195_ ;
  assign \new_Sorter100|17295_  = \new_Sorter100|17194_  | \new_Sorter100|17195_ ;
  assign \new_Sorter100|17296_  = \new_Sorter100|17196_  & \new_Sorter100|17197_ ;
  assign \new_Sorter100|17297_  = \new_Sorter100|17196_  | \new_Sorter100|17197_ ;
  assign \new_Sorter100|17298_  = \new_Sorter100|17198_  & \new_Sorter100|17199_ ;
  assign \new_Sorter100|17299_  = \new_Sorter100|17198_  | \new_Sorter100|17199_ ;
  assign \new_Sorter100|17300_  = \new_Sorter100|17200_ ;
  assign \new_Sorter100|17399_  = \new_Sorter100|17299_ ;
  assign \new_Sorter100|17301_  = \new_Sorter100|17201_  & \new_Sorter100|17202_ ;
  assign \new_Sorter100|17302_  = \new_Sorter100|17201_  | \new_Sorter100|17202_ ;
  assign \new_Sorter100|17303_  = \new_Sorter100|17203_  & \new_Sorter100|17204_ ;
  assign \new_Sorter100|17304_  = \new_Sorter100|17203_  | \new_Sorter100|17204_ ;
  assign \new_Sorter100|17305_  = \new_Sorter100|17205_  & \new_Sorter100|17206_ ;
  assign \new_Sorter100|17306_  = \new_Sorter100|17205_  | \new_Sorter100|17206_ ;
  assign \new_Sorter100|17307_  = \new_Sorter100|17207_  & \new_Sorter100|17208_ ;
  assign \new_Sorter100|17308_  = \new_Sorter100|17207_  | \new_Sorter100|17208_ ;
  assign \new_Sorter100|17309_  = \new_Sorter100|17209_  & \new_Sorter100|17210_ ;
  assign \new_Sorter100|17310_  = \new_Sorter100|17209_  | \new_Sorter100|17210_ ;
  assign \new_Sorter100|17311_  = \new_Sorter100|17211_  & \new_Sorter100|17212_ ;
  assign \new_Sorter100|17312_  = \new_Sorter100|17211_  | \new_Sorter100|17212_ ;
  assign \new_Sorter100|17313_  = \new_Sorter100|17213_  & \new_Sorter100|17214_ ;
  assign \new_Sorter100|17314_  = \new_Sorter100|17213_  | \new_Sorter100|17214_ ;
  assign \new_Sorter100|17315_  = \new_Sorter100|17215_  & \new_Sorter100|17216_ ;
  assign \new_Sorter100|17316_  = \new_Sorter100|17215_  | \new_Sorter100|17216_ ;
  assign \new_Sorter100|17317_  = \new_Sorter100|17217_  & \new_Sorter100|17218_ ;
  assign \new_Sorter100|17318_  = \new_Sorter100|17217_  | \new_Sorter100|17218_ ;
  assign \new_Sorter100|17319_  = \new_Sorter100|17219_  & \new_Sorter100|17220_ ;
  assign \new_Sorter100|17320_  = \new_Sorter100|17219_  | \new_Sorter100|17220_ ;
  assign \new_Sorter100|17321_  = \new_Sorter100|17221_  & \new_Sorter100|17222_ ;
  assign \new_Sorter100|17322_  = \new_Sorter100|17221_  | \new_Sorter100|17222_ ;
  assign \new_Sorter100|17323_  = \new_Sorter100|17223_  & \new_Sorter100|17224_ ;
  assign \new_Sorter100|17324_  = \new_Sorter100|17223_  | \new_Sorter100|17224_ ;
  assign \new_Sorter100|17325_  = \new_Sorter100|17225_  & \new_Sorter100|17226_ ;
  assign \new_Sorter100|17326_  = \new_Sorter100|17225_  | \new_Sorter100|17226_ ;
  assign \new_Sorter100|17327_  = \new_Sorter100|17227_  & \new_Sorter100|17228_ ;
  assign \new_Sorter100|17328_  = \new_Sorter100|17227_  | \new_Sorter100|17228_ ;
  assign \new_Sorter100|17329_  = \new_Sorter100|17229_  & \new_Sorter100|17230_ ;
  assign \new_Sorter100|17330_  = \new_Sorter100|17229_  | \new_Sorter100|17230_ ;
  assign \new_Sorter100|17331_  = \new_Sorter100|17231_  & \new_Sorter100|17232_ ;
  assign \new_Sorter100|17332_  = \new_Sorter100|17231_  | \new_Sorter100|17232_ ;
  assign \new_Sorter100|17333_  = \new_Sorter100|17233_  & \new_Sorter100|17234_ ;
  assign \new_Sorter100|17334_  = \new_Sorter100|17233_  | \new_Sorter100|17234_ ;
  assign \new_Sorter100|17335_  = \new_Sorter100|17235_  & \new_Sorter100|17236_ ;
  assign \new_Sorter100|17336_  = \new_Sorter100|17235_  | \new_Sorter100|17236_ ;
  assign \new_Sorter100|17337_  = \new_Sorter100|17237_  & \new_Sorter100|17238_ ;
  assign \new_Sorter100|17338_  = \new_Sorter100|17237_  | \new_Sorter100|17238_ ;
  assign \new_Sorter100|17339_  = \new_Sorter100|17239_  & \new_Sorter100|17240_ ;
  assign \new_Sorter100|17340_  = \new_Sorter100|17239_  | \new_Sorter100|17240_ ;
  assign \new_Sorter100|17341_  = \new_Sorter100|17241_  & \new_Sorter100|17242_ ;
  assign \new_Sorter100|17342_  = \new_Sorter100|17241_  | \new_Sorter100|17242_ ;
  assign \new_Sorter100|17343_  = \new_Sorter100|17243_  & \new_Sorter100|17244_ ;
  assign \new_Sorter100|17344_  = \new_Sorter100|17243_  | \new_Sorter100|17244_ ;
  assign \new_Sorter100|17345_  = \new_Sorter100|17245_  & \new_Sorter100|17246_ ;
  assign \new_Sorter100|17346_  = \new_Sorter100|17245_  | \new_Sorter100|17246_ ;
  assign \new_Sorter100|17347_  = \new_Sorter100|17247_  & \new_Sorter100|17248_ ;
  assign \new_Sorter100|17348_  = \new_Sorter100|17247_  | \new_Sorter100|17248_ ;
  assign \new_Sorter100|17349_  = \new_Sorter100|17249_  & \new_Sorter100|17250_ ;
  assign \new_Sorter100|17350_  = \new_Sorter100|17249_  | \new_Sorter100|17250_ ;
  assign \new_Sorter100|17351_  = \new_Sorter100|17251_  & \new_Sorter100|17252_ ;
  assign \new_Sorter100|17352_  = \new_Sorter100|17251_  | \new_Sorter100|17252_ ;
  assign \new_Sorter100|17353_  = \new_Sorter100|17253_  & \new_Sorter100|17254_ ;
  assign \new_Sorter100|17354_  = \new_Sorter100|17253_  | \new_Sorter100|17254_ ;
  assign \new_Sorter100|17355_  = \new_Sorter100|17255_  & \new_Sorter100|17256_ ;
  assign \new_Sorter100|17356_  = \new_Sorter100|17255_  | \new_Sorter100|17256_ ;
  assign \new_Sorter100|17357_  = \new_Sorter100|17257_  & \new_Sorter100|17258_ ;
  assign \new_Sorter100|17358_  = \new_Sorter100|17257_  | \new_Sorter100|17258_ ;
  assign \new_Sorter100|17359_  = \new_Sorter100|17259_  & \new_Sorter100|17260_ ;
  assign \new_Sorter100|17360_  = \new_Sorter100|17259_  | \new_Sorter100|17260_ ;
  assign \new_Sorter100|17361_  = \new_Sorter100|17261_  & \new_Sorter100|17262_ ;
  assign \new_Sorter100|17362_  = \new_Sorter100|17261_  | \new_Sorter100|17262_ ;
  assign \new_Sorter100|17363_  = \new_Sorter100|17263_  & \new_Sorter100|17264_ ;
  assign \new_Sorter100|17364_  = \new_Sorter100|17263_  | \new_Sorter100|17264_ ;
  assign \new_Sorter100|17365_  = \new_Sorter100|17265_  & \new_Sorter100|17266_ ;
  assign \new_Sorter100|17366_  = \new_Sorter100|17265_  | \new_Sorter100|17266_ ;
  assign \new_Sorter100|17367_  = \new_Sorter100|17267_  & \new_Sorter100|17268_ ;
  assign \new_Sorter100|17368_  = \new_Sorter100|17267_  | \new_Sorter100|17268_ ;
  assign \new_Sorter100|17369_  = \new_Sorter100|17269_  & \new_Sorter100|17270_ ;
  assign \new_Sorter100|17370_  = \new_Sorter100|17269_  | \new_Sorter100|17270_ ;
  assign \new_Sorter100|17371_  = \new_Sorter100|17271_  & \new_Sorter100|17272_ ;
  assign \new_Sorter100|17372_  = \new_Sorter100|17271_  | \new_Sorter100|17272_ ;
  assign \new_Sorter100|17373_  = \new_Sorter100|17273_  & \new_Sorter100|17274_ ;
  assign \new_Sorter100|17374_  = \new_Sorter100|17273_  | \new_Sorter100|17274_ ;
  assign \new_Sorter100|17375_  = \new_Sorter100|17275_  & \new_Sorter100|17276_ ;
  assign \new_Sorter100|17376_  = \new_Sorter100|17275_  | \new_Sorter100|17276_ ;
  assign \new_Sorter100|17377_  = \new_Sorter100|17277_  & \new_Sorter100|17278_ ;
  assign \new_Sorter100|17378_  = \new_Sorter100|17277_  | \new_Sorter100|17278_ ;
  assign \new_Sorter100|17379_  = \new_Sorter100|17279_  & \new_Sorter100|17280_ ;
  assign \new_Sorter100|17380_  = \new_Sorter100|17279_  | \new_Sorter100|17280_ ;
  assign \new_Sorter100|17381_  = \new_Sorter100|17281_  & \new_Sorter100|17282_ ;
  assign \new_Sorter100|17382_  = \new_Sorter100|17281_  | \new_Sorter100|17282_ ;
  assign \new_Sorter100|17383_  = \new_Sorter100|17283_  & \new_Sorter100|17284_ ;
  assign \new_Sorter100|17384_  = \new_Sorter100|17283_  | \new_Sorter100|17284_ ;
  assign \new_Sorter100|17385_  = \new_Sorter100|17285_  & \new_Sorter100|17286_ ;
  assign \new_Sorter100|17386_  = \new_Sorter100|17285_  | \new_Sorter100|17286_ ;
  assign \new_Sorter100|17387_  = \new_Sorter100|17287_  & \new_Sorter100|17288_ ;
  assign \new_Sorter100|17388_  = \new_Sorter100|17287_  | \new_Sorter100|17288_ ;
  assign \new_Sorter100|17389_  = \new_Sorter100|17289_  & \new_Sorter100|17290_ ;
  assign \new_Sorter100|17390_  = \new_Sorter100|17289_  | \new_Sorter100|17290_ ;
  assign \new_Sorter100|17391_  = \new_Sorter100|17291_  & \new_Sorter100|17292_ ;
  assign \new_Sorter100|17392_  = \new_Sorter100|17291_  | \new_Sorter100|17292_ ;
  assign \new_Sorter100|17393_  = \new_Sorter100|17293_  & \new_Sorter100|17294_ ;
  assign \new_Sorter100|17394_  = \new_Sorter100|17293_  | \new_Sorter100|17294_ ;
  assign \new_Sorter100|17395_  = \new_Sorter100|17295_  & \new_Sorter100|17296_ ;
  assign \new_Sorter100|17396_  = \new_Sorter100|17295_  | \new_Sorter100|17296_ ;
  assign \new_Sorter100|17397_  = \new_Sorter100|17297_  & \new_Sorter100|17298_ ;
  assign \new_Sorter100|17398_  = \new_Sorter100|17297_  | \new_Sorter100|17298_ ;
  assign \new_Sorter100|17400_  = \new_Sorter100|17300_  & \new_Sorter100|17301_ ;
  assign \new_Sorter100|17401_  = \new_Sorter100|17300_  | \new_Sorter100|17301_ ;
  assign \new_Sorter100|17402_  = \new_Sorter100|17302_  & \new_Sorter100|17303_ ;
  assign \new_Sorter100|17403_  = \new_Sorter100|17302_  | \new_Sorter100|17303_ ;
  assign \new_Sorter100|17404_  = \new_Sorter100|17304_  & \new_Sorter100|17305_ ;
  assign \new_Sorter100|17405_  = \new_Sorter100|17304_  | \new_Sorter100|17305_ ;
  assign \new_Sorter100|17406_  = \new_Sorter100|17306_  & \new_Sorter100|17307_ ;
  assign \new_Sorter100|17407_  = \new_Sorter100|17306_  | \new_Sorter100|17307_ ;
  assign \new_Sorter100|17408_  = \new_Sorter100|17308_  & \new_Sorter100|17309_ ;
  assign \new_Sorter100|17409_  = \new_Sorter100|17308_  | \new_Sorter100|17309_ ;
  assign \new_Sorter100|17410_  = \new_Sorter100|17310_  & \new_Sorter100|17311_ ;
  assign \new_Sorter100|17411_  = \new_Sorter100|17310_  | \new_Sorter100|17311_ ;
  assign \new_Sorter100|17412_  = \new_Sorter100|17312_  & \new_Sorter100|17313_ ;
  assign \new_Sorter100|17413_  = \new_Sorter100|17312_  | \new_Sorter100|17313_ ;
  assign \new_Sorter100|17414_  = \new_Sorter100|17314_  & \new_Sorter100|17315_ ;
  assign \new_Sorter100|17415_  = \new_Sorter100|17314_  | \new_Sorter100|17315_ ;
  assign \new_Sorter100|17416_  = \new_Sorter100|17316_  & \new_Sorter100|17317_ ;
  assign \new_Sorter100|17417_  = \new_Sorter100|17316_  | \new_Sorter100|17317_ ;
  assign \new_Sorter100|17418_  = \new_Sorter100|17318_  & \new_Sorter100|17319_ ;
  assign \new_Sorter100|17419_  = \new_Sorter100|17318_  | \new_Sorter100|17319_ ;
  assign \new_Sorter100|17420_  = \new_Sorter100|17320_  & \new_Sorter100|17321_ ;
  assign \new_Sorter100|17421_  = \new_Sorter100|17320_  | \new_Sorter100|17321_ ;
  assign \new_Sorter100|17422_  = \new_Sorter100|17322_  & \new_Sorter100|17323_ ;
  assign \new_Sorter100|17423_  = \new_Sorter100|17322_  | \new_Sorter100|17323_ ;
  assign \new_Sorter100|17424_  = \new_Sorter100|17324_  & \new_Sorter100|17325_ ;
  assign \new_Sorter100|17425_  = \new_Sorter100|17324_  | \new_Sorter100|17325_ ;
  assign \new_Sorter100|17426_  = \new_Sorter100|17326_  & \new_Sorter100|17327_ ;
  assign \new_Sorter100|17427_  = \new_Sorter100|17326_  | \new_Sorter100|17327_ ;
  assign \new_Sorter100|17428_  = \new_Sorter100|17328_  & \new_Sorter100|17329_ ;
  assign \new_Sorter100|17429_  = \new_Sorter100|17328_  | \new_Sorter100|17329_ ;
  assign \new_Sorter100|17430_  = \new_Sorter100|17330_  & \new_Sorter100|17331_ ;
  assign \new_Sorter100|17431_  = \new_Sorter100|17330_  | \new_Sorter100|17331_ ;
  assign \new_Sorter100|17432_  = \new_Sorter100|17332_  & \new_Sorter100|17333_ ;
  assign \new_Sorter100|17433_  = \new_Sorter100|17332_  | \new_Sorter100|17333_ ;
  assign \new_Sorter100|17434_  = \new_Sorter100|17334_  & \new_Sorter100|17335_ ;
  assign \new_Sorter100|17435_  = \new_Sorter100|17334_  | \new_Sorter100|17335_ ;
  assign \new_Sorter100|17436_  = \new_Sorter100|17336_  & \new_Sorter100|17337_ ;
  assign \new_Sorter100|17437_  = \new_Sorter100|17336_  | \new_Sorter100|17337_ ;
  assign \new_Sorter100|17438_  = \new_Sorter100|17338_  & \new_Sorter100|17339_ ;
  assign \new_Sorter100|17439_  = \new_Sorter100|17338_  | \new_Sorter100|17339_ ;
  assign \new_Sorter100|17440_  = \new_Sorter100|17340_  & \new_Sorter100|17341_ ;
  assign \new_Sorter100|17441_  = \new_Sorter100|17340_  | \new_Sorter100|17341_ ;
  assign \new_Sorter100|17442_  = \new_Sorter100|17342_  & \new_Sorter100|17343_ ;
  assign \new_Sorter100|17443_  = \new_Sorter100|17342_  | \new_Sorter100|17343_ ;
  assign \new_Sorter100|17444_  = \new_Sorter100|17344_  & \new_Sorter100|17345_ ;
  assign \new_Sorter100|17445_  = \new_Sorter100|17344_  | \new_Sorter100|17345_ ;
  assign \new_Sorter100|17446_  = \new_Sorter100|17346_  & \new_Sorter100|17347_ ;
  assign \new_Sorter100|17447_  = \new_Sorter100|17346_  | \new_Sorter100|17347_ ;
  assign \new_Sorter100|17448_  = \new_Sorter100|17348_  & \new_Sorter100|17349_ ;
  assign \new_Sorter100|17449_  = \new_Sorter100|17348_  | \new_Sorter100|17349_ ;
  assign \new_Sorter100|17450_  = \new_Sorter100|17350_  & \new_Sorter100|17351_ ;
  assign \new_Sorter100|17451_  = \new_Sorter100|17350_  | \new_Sorter100|17351_ ;
  assign \new_Sorter100|17452_  = \new_Sorter100|17352_  & \new_Sorter100|17353_ ;
  assign \new_Sorter100|17453_  = \new_Sorter100|17352_  | \new_Sorter100|17353_ ;
  assign \new_Sorter100|17454_  = \new_Sorter100|17354_  & \new_Sorter100|17355_ ;
  assign \new_Sorter100|17455_  = \new_Sorter100|17354_  | \new_Sorter100|17355_ ;
  assign \new_Sorter100|17456_  = \new_Sorter100|17356_  & \new_Sorter100|17357_ ;
  assign \new_Sorter100|17457_  = \new_Sorter100|17356_  | \new_Sorter100|17357_ ;
  assign \new_Sorter100|17458_  = \new_Sorter100|17358_  & \new_Sorter100|17359_ ;
  assign \new_Sorter100|17459_  = \new_Sorter100|17358_  | \new_Sorter100|17359_ ;
  assign \new_Sorter100|17460_  = \new_Sorter100|17360_  & \new_Sorter100|17361_ ;
  assign \new_Sorter100|17461_  = \new_Sorter100|17360_  | \new_Sorter100|17361_ ;
  assign \new_Sorter100|17462_  = \new_Sorter100|17362_  & \new_Sorter100|17363_ ;
  assign \new_Sorter100|17463_  = \new_Sorter100|17362_  | \new_Sorter100|17363_ ;
  assign \new_Sorter100|17464_  = \new_Sorter100|17364_  & \new_Sorter100|17365_ ;
  assign \new_Sorter100|17465_  = \new_Sorter100|17364_  | \new_Sorter100|17365_ ;
  assign \new_Sorter100|17466_  = \new_Sorter100|17366_  & \new_Sorter100|17367_ ;
  assign \new_Sorter100|17467_  = \new_Sorter100|17366_  | \new_Sorter100|17367_ ;
  assign \new_Sorter100|17468_  = \new_Sorter100|17368_  & \new_Sorter100|17369_ ;
  assign \new_Sorter100|17469_  = \new_Sorter100|17368_  | \new_Sorter100|17369_ ;
  assign \new_Sorter100|17470_  = \new_Sorter100|17370_  & \new_Sorter100|17371_ ;
  assign \new_Sorter100|17471_  = \new_Sorter100|17370_  | \new_Sorter100|17371_ ;
  assign \new_Sorter100|17472_  = \new_Sorter100|17372_  & \new_Sorter100|17373_ ;
  assign \new_Sorter100|17473_  = \new_Sorter100|17372_  | \new_Sorter100|17373_ ;
  assign \new_Sorter100|17474_  = \new_Sorter100|17374_  & \new_Sorter100|17375_ ;
  assign \new_Sorter100|17475_  = \new_Sorter100|17374_  | \new_Sorter100|17375_ ;
  assign \new_Sorter100|17476_  = \new_Sorter100|17376_  & \new_Sorter100|17377_ ;
  assign \new_Sorter100|17477_  = \new_Sorter100|17376_  | \new_Sorter100|17377_ ;
  assign \new_Sorter100|17478_  = \new_Sorter100|17378_  & \new_Sorter100|17379_ ;
  assign \new_Sorter100|17479_  = \new_Sorter100|17378_  | \new_Sorter100|17379_ ;
  assign \new_Sorter100|17480_  = \new_Sorter100|17380_  & \new_Sorter100|17381_ ;
  assign \new_Sorter100|17481_  = \new_Sorter100|17380_  | \new_Sorter100|17381_ ;
  assign \new_Sorter100|17482_  = \new_Sorter100|17382_  & \new_Sorter100|17383_ ;
  assign \new_Sorter100|17483_  = \new_Sorter100|17382_  | \new_Sorter100|17383_ ;
  assign \new_Sorter100|17484_  = \new_Sorter100|17384_  & \new_Sorter100|17385_ ;
  assign \new_Sorter100|17485_  = \new_Sorter100|17384_  | \new_Sorter100|17385_ ;
  assign \new_Sorter100|17486_  = \new_Sorter100|17386_  & \new_Sorter100|17387_ ;
  assign \new_Sorter100|17487_  = \new_Sorter100|17386_  | \new_Sorter100|17387_ ;
  assign \new_Sorter100|17488_  = \new_Sorter100|17388_  & \new_Sorter100|17389_ ;
  assign \new_Sorter100|17489_  = \new_Sorter100|17388_  | \new_Sorter100|17389_ ;
  assign \new_Sorter100|17490_  = \new_Sorter100|17390_  & \new_Sorter100|17391_ ;
  assign \new_Sorter100|17491_  = \new_Sorter100|17390_  | \new_Sorter100|17391_ ;
  assign \new_Sorter100|17492_  = \new_Sorter100|17392_  & \new_Sorter100|17393_ ;
  assign \new_Sorter100|17493_  = \new_Sorter100|17392_  | \new_Sorter100|17393_ ;
  assign \new_Sorter100|17494_  = \new_Sorter100|17394_  & \new_Sorter100|17395_ ;
  assign \new_Sorter100|17495_  = \new_Sorter100|17394_  | \new_Sorter100|17395_ ;
  assign \new_Sorter100|17496_  = \new_Sorter100|17396_  & \new_Sorter100|17397_ ;
  assign \new_Sorter100|17497_  = \new_Sorter100|17396_  | \new_Sorter100|17397_ ;
  assign \new_Sorter100|17498_  = \new_Sorter100|17398_  & \new_Sorter100|17399_ ;
  assign \new_Sorter100|17499_  = \new_Sorter100|17398_  | \new_Sorter100|17399_ ;
  assign \new_Sorter100|17500_  = \new_Sorter100|17400_ ;
  assign \new_Sorter100|17599_  = \new_Sorter100|17499_ ;
  assign \new_Sorter100|17501_  = \new_Sorter100|17401_  & \new_Sorter100|17402_ ;
  assign \new_Sorter100|17502_  = \new_Sorter100|17401_  | \new_Sorter100|17402_ ;
  assign \new_Sorter100|17503_  = \new_Sorter100|17403_  & \new_Sorter100|17404_ ;
  assign \new_Sorter100|17504_  = \new_Sorter100|17403_  | \new_Sorter100|17404_ ;
  assign \new_Sorter100|17505_  = \new_Sorter100|17405_  & \new_Sorter100|17406_ ;
  assign \new_Sorter100|17506_  = \new_Sorter100|17405_  | \new_Sorter100|17406_ ;
  assign \new_Sorter100|17507_  = \new_Sorter100|17407_  & \new_Sorter100|17408_ ;
  assign \new_Sorter100|17508_  = \new_Sorter100|17407_  | \new_Sorter100|17408_ ;
  assign \new_Sorter100|17509_  = \new_Sorter100|17409_  & \new_Sorter100|17410_ ;
  assign \new_Sorter100|17510_  = \new_Sorter100|17409_  | \new_Sorter100|17410_ ;
  assign \new_Sorter100|17511_  = \new_Sorter100|17411_  & \new_Sorter100|17412_ ;
  assign \new_Sorter100|17512_  = \new_Sorter100|17411_  | \new_Sorter100|17412_ ;
  assign \new_Sorter100|17513_  = \new_Sorter100|17413_  & \new_Sorter100|17414_ ;
  assign \new_Sorter100|17514_  = \new_Sorter100|17413_  | \new_Sorter100|17414_ ;
  assign \new_Sorter100|17515_  = \new_Sorter100|17415_  & \new_Sorter100|17416_ ;
  assign \new_Sorter100|17516_  = \new_Sorter100|17415_  | \new_Sorter100|17416_ ;
  assign \new_Sorter100|17517_  = \new_Sorter100|17417_  & \new_Sorter100|17418_ ;
  assign \new_Sorter100|17518_  = \new_Sorter100|17417_  | \new_Sorter100|17418_ ;
  assign \new_Sorter100|17519_  = \new_Sorter100|17419_  & \new_Sorter100|17420_ ;
  assign \new_Sorter100|17520_  = \new_Sorter100|17419_  | \new_Sorter100|17420_ ;
  assign \new_Sorter100|17521_  = \new_Sorter100|17421_  & \new_Sorter100|17422_ ;
  assign \new_Sorter100|17522_  = \new_Sorter100|17421_  | \new_Sorter100|17422_ ;
  assign \new_Sorter100|17523_  = \new_Sorter100|17423_  & \new_Sorter100|17424_ ;
  assign \new_Sorter100|17524_  = \new_Sorter100|17423_  | \new_Sorter100|17424_ ;
  assign \new_Sorter100|17525_  = \new_Sorter100|17425_  & \new_Sorter100|17426_ ;
  assign \new_Sorter100|17526_  = \new_Sorter100|17425_  | \new_Sorter100|17426_ ;
  assign \new_Sorter100|17527_  = \new_Sorter100|17427_  & \new_Sorter100|17428_ ;
  assign \new_Sorter100|17528_  = \new_Sorter100|17427_  | \new_Sorter100|17428_ ;
  assign \new_Sorter100|17529_  = \new_Sorter100|17429_  & \new_Sorter100|17430_ ;
  assign \new_Sorter100|17530_  = \new_Sorter100|17429_  | \new_Sorter100|17430_ ;
  assign \new_Sorter100|17531_  = \new_Sorter100|17431_  & \new_Sorter100|17432_ ;
  assign \new_Sorter100|17532_  = \new_Sorter100|17431_  | \new_Sorter100|17432_ ;
  assign \new_Sorter100|17533_  = \new_Sorter100|17433_  & \new_Sorter100|17434_ ;
  assign \new_Sorter100|17534_  = \new_Sorter100|17433_  | \new_Sorter100|17434_ ;
  assign \new_Sorter100|17535_  = \new_Sorter100|17435_  & \new_Sorter100|17436_ ;
  assign \new_Sorter100|17536_  = \new_Sorter100|17435_  | \new_Sorter100|17436_ ;
  assign \new_Sorter100|17537_  = \new_Sorter100|17437_  & \new_Sorter100|17438_ ;
  assign \new_Sorter100|17538_  = \new_Sorter100|17437_  | \new_Sorter100|17438_ ;
  assign \new_Sorter100|17539_  = \new_Sorter100|17439_  & \new_Sorter100|17440_ ;
  assign \new_Sorter100|17540_  = \new_Sorter100|17439_  | \new_Sorter100|17440_ ;
  assign \new_Sorter100|17541_  = \new_Sorter100|17441_  & \new_Sorter100|17442_ ;
  assign \new_Sorter100|17542_  = \new_Sorter100|17441_  | \new_Sorter100|17442_ ;
  assign \new_Sorter100|17543_  = \new_Sorter100|17443_  & \new_Sorter100|17444_ ;
  assign \new_Sorter100|17544_  = \new_Sorter100|17443_  | \new_Sorter100|17444_ ;
  assign \new_Sorter100|17545_  = \new_Sorter100|17445_  & \new_Sorter100|17446_ ;
  assign \new_Sorter100|17546_  = \new_Sorter100|17445_  | \new_Sorter100|17446_ ;
  assign \new_Sorter100|17547_  = \new_Sorter100|17447_  & \new_Sorter100|17448_ ;
  assign \new_Sorter100|17548_  = \new_Sorter100|17447_  | \new_Sorter100|17448_ ;
  assign \new_Sorter100|17549_  = \new_Sorter100|17449_  & \new_Sorter100|17450_ ;
  assign \new_Sorter100|17550_  = \new_Sorter100|17449_  | \new_Sorter100|17450_ ;
  assign \new_Sorter100|17551_  = \new_Sorter100|17451_  & \new_Sorter100|17452_ ;
  assign \new_Sorter100|17552_  = \new_Sorter100|17451_  | \new_Sorter100|17452_ ;
  assign \new_Sorter100|17553_  = \new_Sorter100|17453_  & \new_Sorter100|17454_ ;
  assign \new_Sorter100|17554_  = \new_Sorter100|17453_  | \new_Sorter100|17454_ ;
  assign \new_Sorter100|17555_  = \new_Sorter100|17455_  & \new_Sorter100|17456_ ;
  assign \new_Sorter100|17556_  = \new_Sorter100|17455_  | \new_Sorter100|17456_ ;
  assign \new_Sorter100|17557_  = \new_Sorter100|17457_  & \new_Sorter100|17458_ ;
  assign \new_Sorter100|17558_  = \new_Sorter100|17457_  | \new_Sorter100|17458_ ;
  assign \new_Sorter100|17559_  = \new_Sorter100|17459_  & \new_Sorter100|17460_ ;
  assign \new_Sorter100|17560_  = \new_Sorter100|17459_  | \new_Sorter100|17460_ ;
  assign \new_Sorter100|17561_  = \new_Sorter100|17461_  & \new_Sorter100|17462_ ;
  assign \new_Sorter100|17562_  = \new_Sorter100|17461_  | \new_Sorter100|17462_ ;
  assign \new_Sorter100|17563_  = \new_Sorter100|17463_  & \new_Sorter100|17464_ ;
  assign \new_Sorter100|17564_  = \new_Sorter100|17463_  | \new_Sorter100|17464_ ;
  assign \new_Sorter100|17565_  = \new_Sorter100|17465_  & \new_Sorter100|17466_ ;
  assign \new_Sorter100|17566_  = \new_Sorter100|17465_  | \new_Sorter100|17466_ ;
  assign \new_Sorter100|17567_  = \new_Sorter100|17467_  & \new_Sorter100|17468_ ;
  assign \new_Sorter100|17568_  = \new_Sorter100|17467_  | \new_Sorter100|17468_ ;
  assign \new_Sorter100|17569_  = \new_Sorter100|17469_  & \new_Sorter100|17470_ ;
  assign \new_Sorter100|17570_  = \new_Sorter100|17469_  | \new_Sorter100|17470_ ;
  assign \new_Sorter100|17571_  = \new_Sorter100|17471_  & \new_Sorter100|17472_ ;
  assign \new_Sorter100|17572_  = \new_Sorter100|17471_  | \new_Sorter100|17472_ ;
  assign \new_Sorter100|17573_  = \new_Sorter100|17473_  & \new_Sorter100|17474_ ;
  assign \new_Sorter100|17574_  = \new_Sorter100|17473_  | \new_Sorter100|17474_ ;
  assign \new_Sorter100|17575_  = \new_Sorter100|17475_  & \new_Sorter100|17476_ ;
  assign \new_Sorter100|17576_  = \new_Sorter100|17475_  | \new_Sorter100|17476_ ;
  assign \new_Sorter100|17577_  = \new_Sorter100|17477_  & \new_Sorter100|17478_ ;
  assign \new_Sorter100|17578_  = \new_Sorter100|17477_  | \new_Sorter100|17478_ ;
  assign \new_Sorter100|17579_  = \new_Sorter100|17479_  & \new_Sorter100|17480_ ;
  assign \new_Sorter100|17580_  = \new_Sorter100|17479_  | \new_Sorter100|17480_ ;
  assign \new_Sorter100|17581_  = \new_Sorter100|17481_  & \new_Sorter100|17482_ ;
  assign \new_Sorter100|17582_  = \new_Sorter100|17481_  | \new_Sorter100|17482_ ;
  assign \new_Sorter100|17583_  = \new_Sorter100|17483_  & \new_Sorter100|17484_ ;
  assign \new_Sorter100|17584_  = \new_Sorter100|17483_  | \new_Sorter100|17484_ ;
  assign \new_Sorter100|17585_  = \new_Sorter100|17485_  & \new_Sorter100|17486_ ;
  assign \new_Sorter100|17586_  = \new_Sorter100|17485_  | \new_Sorter100|17486_ ;
  assign \new_Sorter100|17587_  = \new_Sorter100|17487_  & \new_Sorter100|17488_ ;
  assign \new_Sorter100|17588_  = \new_Sorter100|17487_  | \new_Sorter100|17488_ ;
  assign \new_Sorter100|17589_  = \new_Sorter100|17489_  & \new_Sorter100|17490_ ;
  assign \new_Sorter100|17590_  = \new_Sorter100|17489_  | \new_Sorter100|17490_ ;
  assign \new_Sorter100|17591_  = \new_Sorter100|17491_  & \new_Sorter100|17492_ ;
  assign \new_Sorter100|17592_  = \new_Sorter100|17491_  | \new_Sorter100|17492_ ;
  assign \new_Sorter100|17593_  = \new_Sorter100|17493_  & \new_Sorter100|17494_ ;
  assign \new_Sorter100|17594_  = \new_Sorter100|17493_  | \new_Sorter100|17494_ ;
  assign \new_Sorter100|17595_  = \new_Sorter100|17495_  & \new_Sorter100|17496_ ;
  assign \new_Sorter100|17596_  = \new_Sorter100|17495_  | \new_Sorter100|17496_ ;
  assign \new_Sorter100|17597_  = \new_Sorter100|17497_  & \new_Sorter100|17498_ ;
  assign \new_Sorter100|17598_  = \new_Sorter100|17497_  | \new_Sorter100|17498_ ;
  assign \new_Sorter100|17600_  = \new_Sorter100|17500_  & \new_Sorter100|17501_ ;
  assign \new_Sorter100|17601_  = \new_Sorter100|17500_  | \new_Sorter100|17501_ ;
  assign \new_Sorter100|17602_  = \new_Sorter100|17502_  & \new_Sorter100|17503_ ;
  assign \new_Sorter100|17603_  = \new_Sorter100|17502_  | \new_Sorter100|17503_ ;
  assign \new_Sorter100|17604_  = \new_Sorter100|17504_  & \new_Sorter100|17505_ ;
  assign \new_Sorter100|17605_  = \new_Sorter100|17504_  | \new_Sorter100|17505_ ;
  assign \new_Sorter100|17606_  = \new_Sorter100|17506_  & \new_Sorter100|17507_ ;
  assign \new_Sorter100|17607_  = \new_Sorter100|17506_  | \new_Sorter100|17507_ ;
  assign \new_Sorter100|17608_  = \new_Sorter100|17508_  & \new_Sorter100|17509_ ;
  assign \new_Sorter100|17609_  = \new_Sorter100|17508_  | \new_Sorter100|17509_ ;
  assign \new_Sorter100|17610_  = \new_Sorter100|17510_  & \new_Sorter100|17511_ ;
  assign \new_Sorter100|17611_  = \new_Sorter100|17510_  | \new_Sorter100|17511_ ;
  assign \new_Sorter100|17612_  = \new_Sorter100|17512_  & \new_Sorter100|17513_ ;
  assign \new_Sorter100|17613_  = \new_Sorter100|17512_  | \new_Sorter100|17513_ ;
  assign \new_Sorter100|17614_  = \new_Sorter100|17514_  & \new_Sorter100|17515_ ;
  assign \new_Sorter100|17615_  = \new_Sorter100|17514_  | \new_Sorter100|17515_ ;
  assign \new_Sorter100|17616_  = \new_Sorter100|17516_  & \new_Sorter100|17517_ ;
  assign \new_Sorter100|17617_  = \new_Sorter100|17516_  | \new_Sorter100|17517_ ;
  assign \new_Sorter100|17618_  = \new_Sorter100|17518_  & \new_Sorter100|17519_ ;
  assign \new_Sorter100|17619_  = \new_Sorter100|17518_  | \new_Sorter100|17519_ ;
  assign \new_Sorter100|17620_  = \new_Sorter100|17520_  & \new_Sorter100|17521_ ;
  assign \new_Sorter100|17621_  = \new_Sorter100|17520_  | \new_Sorter100|17521_ ;
  assign \new_Sorter100|17622_  = \new_Sorter100|17522_  & \new_Sorter100|17523_ ;
  assign \new_Sorter100|17623_  = \new_Sorter100|17522_  | \new_Sorter100|17523_ ;
  assign \new_Sorter100|17624_  = \new_Sorter100|17524_  & \new_Sorter100|17525_ ;
  assign \new_Sorter100|17625_  = \new_Sorter100|17524_  | \new_Sorter100|17525_ ;
  assign \new_Sorter100|17626_  = \new_Sorter100|17526_  & \new_Sorter100|17527_ ;
  assign \new_Sorter100|17627_  = \new_Sorter100|17526_  | \new_Sorter100|17527_ ;
  assign \new_Sorter100|17628_  = \new_Sorter100|17528_  & \new_Sorter100|17529_ ;
  assign \new_Sorter100|17629_  = \new_Sorter100|17528_  | \new_Sorter100|17529_ ;
  assign \new_Sorter100|17630_  = \new_Sorter100|17530_  & \new_Sorter100|17531_ ;
  assign \new_Sorter100|17631_  = \new_Sorter100|17530_  | \new_Sorter100|17531_ ;
  assign \new_Sorter100|17632_  = \new_Sorter100|17532_  & \new_Sorter100|17533_ ;
  assign \new_Sorter100|17633_  = \new_Sorter100|17532_  | \new_Sorter100|17533_ ;
  assign \new_Sorter100|17634_  = \new_Sorter100|17534_  & \new_Sorter100|17535_ ;
  assign \new_Sorter100|17635_  = \new_Sorter100|17534_  | \new_Sorter100|17535_ ;
  assign \new_Sorter100|17636_  = \new_Sorter100|17536_  & \new_Sorter100|17537_ ;
  assign \new_Sorter100|17637_  = \new_Sorter100|17536_  | \new_Sorter100|17537_ ;
  assign \new_Sorter100|17638_  = \new_Sorter100|17538_  & \new_Sorter100|17539_ ;
  assign \new_Sorter100|17639_  = \new_Sorter100|17538_  | \new_Sorter100|17539_ ;
  assign \new_Sorter100|17640_  = \new_Sorter100|17540_  & \new_Sorter100|17541_ ;
  assign \new_Sorter100|17641_  = \new_Sorter100|17540_  | \new_Sorter100|17541_ ;
  assign \new_Sorter100|17642_  = \new_Sorter100|17542_  & \new_Sorter100|17543_ ;
  assign \new_Sorter100|17643_  = \new_Sorter100|17542_  | \new_Sorter100|17543_ ;
  assign \new_Sorter100|17644_  = \new_Sorter100|17544_  & \new_Sorter100|17545_ ;
  assign \new_Sorter100|17645_  = \new_Sorter100|17544_  | \new_Sorter100|17545_ ;
  assign \new_Sorter100|17646_  = \new_Sorter100|17546_  & \new_Sorter100|17547_ ;
  assign \new_Sorter100|17647_  = \new_Sorter100|17546_  | \new_Sorter100|17547_ ;
  assign \new_Sorter100|17648_  = \new_Sorter100|17548_  & \new_Sorter100|17549_ ;
  assign \new_Sorter100|17649_  = \new_Sorter100|17548_  | \new_Sorter100|17549_ ;
  assign \new_Sorter100|17650_  = \new_Sorter100|17550_  & \new_Sorter100|17551_ ;
  assign \new_Sorter100|17651_  = \new_Sorter100|17550_  | \new_Sorter100|17551_ ;
  assign \new_Sorter100|17652_  = \new_Sorter100|17552_  & \new_Sorter100|17553_ ;
  assign \new_Sorter100|17653_  = \new_Sorter100|17552_  | \new_Sorter100|17553_ ;
  assign \new_Sorter100|17654_  = \new_Sorter100|17554_  & \new_Sorter100|17555_ ;
  assign \new_Sorter100|17655_  = \new_Sorter100|17554_  | \new_Sorter100|17555_ ;
  assign \new_Sorter100|17656_  = \new_Sorter100|17556_  & \new_Sorter100|17557_ ;
  assign \new_Sorter100|17657_  = \new_Sorter100|17556_  | \new_Sorter100|17557_ ;
  assign \new_Sorter100|17658_  = \new_Sorter100|17558_  & \new_Sorter100|17559_ ;
  assign \new_Sorter100|17659_  = \new_Sorter100|17558_  | \new_Sorter100|17559_ ;
  assign \new_Sorter100|17660_  = \new_Sorter100|17560_  & \new_Sorter100|17561_ ;
  assign \new_Sorter100|17661_  = \new_Sorter100|17560_  | \new_Sorter100|17561_ ;
  assign \new_Sorter100|17662_  = \new_Sorter100|17562_  & \new_Sorter100|17563_ ;
  assign \new_Sorter100|17663_  = \new_Sorter100|17562_  | \new_Sorter100|17563_ ;
  assign \new_Sorter100|17664_  = \new_Sorter100|17564_  & \new_Sorter100|17565_ ;
  assign \new_Sorter100|17665_  = \new_Sorter100|17564_  | \new_Sorter100|17565_ ;
  assign \new_Sorter100|17666_  = \new_Sorter100|17566_  & \new_Sorter100|17567_ ;
  assign \new_Sorter100|17667_  = \new_Sorter100|17566_  | \new_Sorter100|17567_ ;
  assign \new_Sorter100|17668_  = \new_Sorter100|17568_  & \new_Sorter100|17569_ ;
  assign \new_Sorter100|17669_  = \new_Sorter100|17568_  | \new_Sorter100|17569_ ;
  assign \new_Sorter100|17670_  = \new_Sorter100|17570_  & \new_Sorter100|17571_ ;
  assign \new_Sorter100|17671_  = \new_Sorter100|17570_  | \new_Sorter100|17571_ ;
  assign \new_Sorter100|17672_  = \new_Sorter100|17572_  & \new_Sorter100|17573_ ;
  assign \new_Sorter100|17673_  = \new_Sorter100|17572_  | \new_Sorter100|17573_ ;
  assign \new_Sorter100|17674_  = \new_Sorter100|17574_  & \new_Sorter100|17575_ ;
  assign \new_Sorter100|17675_  = \new_Sorter100|17574_  | \new_Sorter100|17575_ ;
  assign \new_Sorter100|17676_  = \new_Sorter100|17576_  & \new_Sorter100|17577_ ;
  assign \new_Sorter100|17677_  = \new_Sorter100|17576_  | \new_Sorter100|17577_ ;
  assign \new_Sorter100|17678_  = \new_Sorter100|17578_  & \new_Sorter100|17579_ ;
  assign \new_Sorter100|17679_  = \new_Sorter100|17578_  | \new_Sorter100|17579_ ;
  assign \new_Sorter100|17680_  = \new_Sorter100|17580_  & \new_Sorter100|17581_ ;
  assign \new_Sorter100|17681_  = \new_Sorter100|17580_  | \new_Sorter100|17581_ ;
  assign \new_Sorter100|17682_  = \new_Sorter100|17582_  & \new_Sorter100|17583_ ;
  assign \new_Sorter100|17683_  = \new_Sorter100|17582_  | \new_Sorter100|17583_ ;
  assign \new_Sorter100|17684_  = \new_Sorter100|17584_  & \new_Sorter100|17585_ ;
  assign \new_Sorter100|17685_  = \new_Sorter100|17584_  | \new_Sorter100|17585_ ;
  assign \new_Sorter100|17686_  = \new_Sorter100|17586_  & \new_Sorter100|17587_ ;
  assign \new_Sorter100|17687_  = \new_Sorter100|17586_  | \new_Sorter100|17587_ ;
  assign \new_Sorter100|17688_  = \new_Sorter100|17588_  & \new_Sorter100|17589_ ;
  assign \new_Sorter100|17689_  = \new_Sorter100|17588_  | \new_Sorter100|17589_ ;
  assign \new_Sorter100|17690_  = \new_Sorter100|17590_  & \new_Sorter100|17591_ ;
  assign \new_Sorter100|17691_  = \new_Sorter100|17590_  | \new_Sorter100|17591_ ;
  assign \new_Sorter100|17692_  = \new_Sorter100|17592_  & \new_Sorter100|17593_ ;
  assign \new_Sorter100|17693_  = \new_Sorter100|17592_  | \new_Sorter100|17593_ ;
  assign \new_Sorter100|17694_  = \new_Sorter100|17594_  & \new_Sorter100|17595_ ;
  assign \new_Sorter100|17695_  = \new_Sorter100|17594_  | \new_Sorter100|17595_ ;
  assign \new_Sorter100|17696_  = \new_Sorter100|17596_  & \new_Sorter100|17597_ ;
  assign \new_Sorter100|17697_  = \new_Sorter100|17596_  | \new_Sorter100|17597_ ;
  assign \new_Sorter100|17698_  = \new_Sorter100|17598_  & \new_Sorter100|17599_ ;
  assign \new_Sorter100|17699_  = \new_Sorter100|17598_  | \new_Sorter100|17599_ ;
  assign \new_Sorter100|17700_  = \new_Sorter100|17600_ ;
  assign \new_Sorter100|17799_  = \new_Sorter100|17699_ ;
  assign \new_Sorter100|17701_  = \new_Sorter100|17601_  & \new_Sorter100|17602_ ;
  assign \new_Sorter100|17702_  = \new_Sorter100|17601_  | \new_Sorter100|17602_ ;
  assign \new_Sorter100|17703_  = \new_Sorter100|17603_  & \new_Sorter100|17604_ ;
  assign \new_Sorter100|17704_  = \new_Sorter100|17603_  | \new_Sorter100|17604_ ;
  assign \new_Sorter100|17705_  = \new_Sorter100|17605_  & \new_Sorter100|17606_ ;
  assign \new_Sorter100|17706_  = \new_Sorter100|17605_  | \new_Sorter100|17606_ ;
  assign \new_Sorter100|17707_  = \new_Sorter100|17607_  & \new_Sorter100|17608_ ;
  assign \new_Sorter100|17708_  = \new_Sorter100|17607_  | \new_Sorter100|17608_ ;
  assign \new_Sorter100|17709_  = \new_Sorter100|17609_  & \new_Sorter100|17610_ ;
  assign \new_Sorter100|17710_  = \new_Sorter100|17609_  | \new_Sorter100|17610_ ;
  assign \new_Sorter100|17711_  = \new_Sorter100|17611_  & \new_Sorter100|17612_ ;
  assign \new_Sorter100|17712_  = \new_Sorter100|17611_  | \new_Sorter100|17612_ ;
  assign \new_Sorter100|17713_  = \new_Sorter100|17613_  & \new_Sorter100|17614_ ;
  assign \new_Sorter100|17714_  = \new_Sorter100|17613_  | \new_Sorter100|17614_ ;
  assign \new_Sorter100|17715_  = \new_Sorter100|17615_  & \new_Sorter100|17616_ ;
  assign \new_Sorter100|17716_  = \new_Sorter100|17615_  | \new_Sorter100|17616_ ;
  assign \new_Sorter100|17717_  = \new_Sorter100|17617_  & \new_Sorter100|17618_ ;
  assign \new_Sorter100|17718_  = \new_Sorter100|17617_  | \new_Sorter100|17618_ ;
  assign \new_Sorter100|17719_  = \new_Sorter100|17619_  & \new_Sorter100|17620_ ;
  assign \new_Sorter100|17720_  = \new_Sorter100|17619_  | \new_Sorter100|17620_ ;
  assign \new_Sorter100|17721_  = \new_Sorter100|17621_  & \new_Sorter100|17622_ ;
  assign \new_Sorter100|17722_  = \new_Sorter100|17621_  | \new_Sorter100|17622_ ;
  assign \new_Sorter100|17723_  = \new_Sorter100|17623_  & \new_Sorter100|17624_ ;
  assign \new_Sorter100|17724_  = \new_Sorter100|17623_  | \new_Sorter100|17624_ ;
  assign \new_Sorter100|17725_  = \new_Sorter100|17625_  & \new_Sorter100|17626_ ;
  assign \new_Sorter100|17726_  = \new_Sorter100|17625_  | \new_Sorter100|17626_ ;
  assign \new_Sorter100|17727_  = \new_Sorter100|17627_  & \new_Sorter100|17628_ ;
  assign \new_Sorter100|17728_  = \new_Sorter100|17627_  | \new_Sorter100|17628_ ;
  assign \new_Sorter100|17729_  = \new_Sorter100|17629_  & \new_Sorter100|17630_ ;
  assign \new_Sorter100|17730_  = \new_Sorter100|17629_  | \new_Sorter100|17630_ ;
  assign \new_Sorter100|17731_  = \new_Sorter100|17631_  & \new_Sorter100|17632_ ;
  assign \new_Sorter100|17732_  = \new_Sorter100|17631_  | \new_Sorter100|17632_ ;
  assign \new_Sorter100|17733_  = \new_Sorter100|17633_  & \new_Sorter100|17634_ ;
  assign \new_Sorter100|17734_  = \new_Sorter100|17633_  | \new_Sorter100|17634_ ;
  assign \new_Sorter100|17735_  = \new_Sorter100|17635_  & \new_Sorter100|17636_ ;
  assign \new_Sorter100|17736_  = \new_Sorter100|17635_  | \new_Sorter100|17636_ ;
  assign \new_Sorter100|17737_  = \new_Sorter100|17637_  & \new_Sorter100|17638_ ;
  assign \new_Sorter100|17738_  = \new_Sorter100|17637_  | \new_Sorter100|17638_ ;
  assign \new_Sorter100|17739_  = \new_Sorter100|17639_  & \new_Sorter100|17640_ ;
  assign \new_Sorter100|17740_  = \new_Sorter100|17639_  | \new_Sorter100|17640_ ;
  assign \new_Sorter100|17741_  = \new_Sorter100|17641_  & \new_Sorter100|17642_ ;
  assign \new_Sorter100|17742_  = \new_Sorter100|17641_  | \new_Sorter100|17642_ ;
  assign \new_Sorter100|17743_  = \new_Sorter100|17643_  & \new_Sorter100|17644_ ;
  assign \new_Sorter100|17744_  = \new_Sorter100|17643_  | \new_Sorter100|17644_ ;
  assign \new_Sorter100|17745_  = \new_Sorter100|17645_  & \new_Sorter100|17646_ ;
  assign \new_Sorter100|17746_  = \new_Sorter100|17645_  | \new_Sorter100|17646_ ;
  assign \new_Sorter100|17747_  = \new_Sorter100|17647_  & \new_Sorter100|17648_ ;
  assign \new_Sorter100|17748_  = \new_Sorter100|17647_  | \new_Sorter100|17648_ ;
  assign \new_Sorter100|17749_  = \new_Sorter100|17649_  & \new_Sorter100|17650_ ;
  assign \new_Sorter100|17750_  = \new_Sorter100|17649_  | \new_Sorter100|17650_ ;
  assign \new_Sorter100|17751_  = \new_Sorter100|17651_  & \new_Sorter100|17652_ ;
  assign \new_Sorter100|17752_  = \new_Sorter100|17651_  | \new_Sorter100|17652_ ;
  assign \new_Sorter100|17753_  = \new_Sorter100|17653_  & \new_Sorter100|17654_ ;
  assign \new_Sorter100|17754_  = \new_Sorter100|17653_  | \new_Sorter100|17654_ ;
  assign \new_Sorter100|17755_  = \new_Sorter100|17655_  & \new_Sorter100|17656_ ;
  assign \new_Sorter100|17756_  = \new_Sorter100|17655_  | \new_Sorter100|17656_ ;
  assign \new_Sorter100|17757_  = \new_Sorter100|17657_  & \new_Sorter100|17658_ ;
  assign \new_Sorter100|17758_  = \new_Sorter100|17657_  | \new_Sorter100|17658_ ;
  assign \new_Sorter100|17759_  = \new_Sorter100|17659_  & \new_Sorter100|17660_ ;
  assign \new_Sorter100|17760_  = \new_Sorter100|17659_  | \new_Sorter100|17660_ ;
  assign \new_Sorter100|17761_  = \new_Sorter100|17661_  & \new_Sorter100|17662_ ;
  assign \new_Sorter100|17762_  = \new_Sorter100|17661_  | \new_Sorter100|17662_ ;
  assign \new_Sorter100|17763_  = \new_Sorter100|17663_  & \new_Sorter100|17664_ ;
  assign \new_Sorter100|17764_  = \new_Sorter100|17663_  | \new_Sorter100|17664_ ;
  assign \new_Sorter100|17765_  = \new_Sorter100|17665_  & \new_Sorter100|17666_ ;
  assign \new_Sorter100|17766_  = \new_Sorter100|17665_  | \new_Sorter100|17666_ ;
  assign \new_Sorter100|17767_  = \new_Sorter100|17667_  & \new_Sorter100|17668_ ;
  assign \new_Sorter100|17768_  = \new_Sorter100|17667_  | \new_Sorter100|17668_ ;
  assign \new_Sorter100|17769_  = \new_Sorter100|17669_  & \new_Sorter100|17670_ ;
  assign \new_Sorter100|17770_  = \new_Sorter100|17669_  | \new_Sorter100|17670_ ;
  assign \new_Sorter100|17771_  = \new_Sorter100|17671_  & \new_Sorter100|17672_ ;
  assign \new_Sorter100|17772_  = \new_Sorter100|17671_  | \new_Sorter100|17672_ ;
  assign \new_Sorter100|17773_  = \new_Sorter100|17673_  & \new_Sorter100|17674_ ;
  assign \new_Sorter100|17774_  = \new_Sorter100|17673_  | \new_Sorter100|17674_ ;
  assign \new_Sorter100|17775_  = \new_Sorter100|17675_  & \new_Sorter100|17676_ ;
  assign \new_Sorter100|17776_  = \new_Sorter100|17675_  | \new_Sorter100|17676_ ;
  assign \new_Sorter100|17777_  = \new_Sorter100|17677_  & \new_Sorter100|17678_ ;
  assign \new_Sorter100|17778_  = \new_Sorter100|17677_  | \new_Sorter100|17678_ ;
  assign \new_Sorter100|17779_  = \new_Sorter100|17679_  & \new_Sorter100|17680_ ;
  assign \new_Sorter100|17780_  = \new_Sorter100|17679_  | \new_Sorter100|17680_ ;
  assign \new_Sorter100|17781_  = \new_Sorter100|17681_  & \new_Sorter100|17682_ ;
  assign \new_Sorter100|17782_  = \new_Sorter100|17681_  | \new_Sorter100|17682_ ;
  assign \new_Sorter100|17783_  = \new_Sorter100|17683_  & \new_Sorter100|17684_ ;
  assign \new_Sorter100|17784_  = \new_Sorter100|17683_  | \new_Sorter100|17684_ ;
  assign \new_Sorter100|17785_  = \new_Sorter100|17685_  & \new_Sorter100|17686_ ;
  assign \new_Sorter100|17786_  = \new_Sorter100|17685_  | \new_Sorter100|17686_ ;
  assign \new_Sorter100|17787_  = \new_Sorter100|17687_  & \new_Sorter100|17688_ ;
  assign \new_Sorter100|17788_  = \new_Sorter100|17687_  | \new_Sorter100|17688_ ;
  assign \new_Sorter100|17789_  = \new_Sorter100|17689_  & \new_Sorter100|17690_ ;
  assign \new_Sorter100|17790_  = \new_Sorter100|17689_  | \new_Sorter100|17690_ ;
  assign \new_Sorter100|17791_  = \new_Sorter100|17691_  & \new_Sorter100|17692_ ;
  assign \new_Sorter100|17792_  = \new_Sorter100|17691_  | \new_Sorter100|17692_ ;
  assign \new_Sorter100|17793_  = \new_Sorter100|17693_  & \new_Sorter100|17694_ ;
  assign \new_Sorter100|17794_  = \new_Sorter100|17693_  | \new_Sorter100|17694_ ;
  assign \new_Sorter100|17795_  = \new_Sorter100|17695_  & \new_Sorter100|17696_ ;
  assign \new_Sorter100|17796_  = \new_Sorter100|17695_  | \new_Sorter100|17696_ ;
  assign \new_Sorter100|17797_  = \new_Sorter100|17697_  & \new_Sorter100|17698_ ;
  assign \new_Sorter100|17798_  = \new_Sorter100|17697_  | \new_Sorter100|17698_ ;
  assign \new_Sorter100|17800_  = \new_Sorter100|17700_  & \new_Sorter100|17701_ ;
  assign \new_Sorter100|17801_  = \new_Sorter100|17700_  | \new_Sorter100|17701_ ;
  assign \new_Sorter100|17802_  = \new_Sorter100|17702_  & \new_Sorter100|17703_ ;
  assign \new_Sorter100|17803_  = \new_Sorter100|17702_  | \new_Sorter100|17703_ ;
  assign \new_Sorter100|17804_  = \new_Sorter100|17704_  & \new_Sorter100|17705_ ;
  assign \new_Sorter100|17805_  = \new_Sorter100|17704_  | \new_Sorter100|17705_ ;
  assign \new_Sorter100|17806_  = \new_Sorter100|17706_  & \new_Sorter100|17707_ ;
  assign \new_Sorter100|17807_  = \new_Sorter100|17706_  | \new_Sorter100|17707_ ;
  assign \new_Sorter100|17808_  = \new_Sorter100|17708_  & \new_Sorter100|17709_ ;
  assign \new_Sorter100|17809_  = \new_Sorter100|17708_  | \new_Sorter100|17709_ ;
  assign \new_Sorter100|17810_  = \new_Sorter100|17710_  & \new_Sorter100|17711_ ;
  assign \new_Sorter100|17811_  = \new_Sorter100|17710_  | \new_Sorter100|17711_ ;
  assign \new_Sorter100|17812_  = \new_Sorter100|17712_  & \new_Sorter100|17713_ ;
  assign \new_Sorter100|17813_  = \new_Sorter100|17712_  | \new_Sorter100|17713_ ;
  assign \new_Sorter100|17814_  = \new_Sorter100|17714_  & \new_Sorter100|17715_ ;
  assign \new_Sorter100|17815_  = \new_Sorter100|17714_  | \new_Sorter100|17715_ ;
  assign \new_Sorter100|17816_  = \new_Sorter100|17716_  & \new_Sorter100|17717_ ;
  assign \new_Sorter100|17817_  = \new_Sorter100|17716_  | \new_Sorter100|17717_ ;
  assign \new_Sorter100|17818_  = \new_Sorter100|17718_  & \new_Sorter100|17719_ ;
  assign \new_Sorter100|17819_  = \new_Sorter100|17718_  | \new_Sorter100|17719_ ;
  assign \new_Sorter100|17820_  = \new_Sorter100|17720_  & \new_Sorter100|17721_ ;
  assign \new_Sorter100|17821_  = \new_Sorter100|17720_  | \new_Sorter100|17721_ ;
  assign \new_Sorter100|17822_  = \new_Sorter100|17722_  & \new_Sorter100|17723_ ;
  assign \new_Sorter100|17823_  = \new_Sorter100|17722_  | \new_Sorter100|17723_ ;
  assign \new_Sorter100|17824_  = \new_Sorter100|17724_  & \new_Sorter100|17725_ ;
  assign \new_Sorter100|17825_  = \new_Sorter100|17724_  | \new_Sorter100|17725_ ;
  assign \new_Sorter100|17826_  = \new_Sorter100|17726_  & \new_Sorter100|17727_ ;
  assign \new_Sorter100|17827_  = \new_Sorter100|17726_  | \new_Sorter100|17727_ ;
  assign \new_Sorter100|17828_  = \new_Sorter100|17728_  & \new_Sorter100|17729_ ;
  assign \new_Sorter100|17829_  = \new_Sorter100|17728_  | \new_Sorter100|17729_ ;
  assign \new_Sorter100|17830_  = \new_Sorter100|17730_  & \new_Sorter100|17731_ ;
  assign \new_Sorter100|17831_  = \new_Sorter100|17730_  | \new_Sorter100|17731_ ;
  assign \new_Sorter100|17832_  = \new_Sorter100|17732_  & \new_Sorter100|17733_ ;
  assign \new_Sorter100|17833_  = \new_Sorter100|17732_  | \new_Sorter100|17733_ ;
  assign \new_Sorter100|17834_  = \new_Sorter100|17734_  & \new_Sorter100|17735_ ;
  assign \new_Sorter100|17835_  = \new_Sorter100|17734_  | \new_Sorter100|17735_ ;
  assign \new_Sorter100|17836_  = \new_Sorter100|17736_  & \new_Sorter100|17737_ ;
  assign \new_Sorter100|17837_  = \new_Sorter100|17736_  | \new_Sorter100|17737_ ;
  assign \new_Sorter100|17838_  = \new_Sorter100|17738_  & \new_Sorter100|17739_ ;
  assign \new_Sorter100|17839_  = \new_Sorter100|17738_  | \new_Sorter100|17739_ ;
  assign \new_Sorter100|17840_  = \new_Sorter100|17740_  & \new_Sorter100|17741_ ;
  assign \new_Sorter100|17841_  = \new_Sorter100|17740_  | \new_Sorter100|17741_ ;
  assign \new_Sorter100|17842_  = \new_Sorter100|17742_  & \new_Sorter100|17743_ ;
  assign \new_Sorter100|17843_  = \new_Sorter100|17742_  | \new_Sorter100|17743_ ;
  assign \new_Sorter100|17844_  = \new_Sorter100|17744_  & \new_Sorter100|17745_ ;
  assign \new_Sorter100|17845_  = \new_Sorter100|17744_  | \new_Sorter100|17745_ ;
  assign \new_Sorter100|17846_  = \new_Sorter100|17746_  & \new_Sorter100|17747_ ;
  assign \new_Sorter100|17847_  = \new_Sorter100|17746_  | \new_Sorter100|17747_ ;
  assign \new_Sorter100|17848_  = \new_Sorter100|17748_  & \new_Sorter100|17749_ ;
  assign \new_Sorter100|17849_  = \new_Sorter100|17748_  | \new_Sorter100|17749_ ;
  assign \new_Sorter100|17850_  = \new_Sorter100|17750_  & \new_Sorter100|17751_ ;
  assign \new_Sorter100|17851_  = \new_Sorter100|17750_  | \new_Sorter100|17751_ ;
  assign \new_Sorter100|17852_  = \new_Sorter100|17752_  & \new_Sorter100|17753_ ;
  assign \new_Sorter100|17853_  = \new_Sorter100|17752_  | \new_Sorter100|17753_ ;
  assign \new_Sorter100|17854_  = \new_Sorter100|17754_  & \new_Sorter100|17755_ ;
  assign \new_Sorter100|17855_  = \new_Sorter100|17754_  | \new_Sorter100|17755_ ;
  assign \new_Sorter100|17856_  = \new_Sorter100|17756_  & \new_Sorter100|17757_ ;
  assign \new_Sorter100|17857_  = \new_Sorter100|17756_  | \new_Sorter100|17757_ ;
  assign \new_Sorter100|17858_  = \new_Sorter100|17758_  & \new_Sorter100|17759_ ;
  assign \new_Sorter100|17859_  = \new_Sorter100|17758_  | \new_Sorter100|17759_ ;
  assign \new_Sorter100|17860_  = \new_Sorter100|17760_  & \new_Sorter100|17761_ ;
  assign \new_Sorter100|17861_  = \new_Sorter100|17760_  | \new_Sorter100|17761_ ;
  assign \new_Sorter100|17862_  = \new_Sorter100|17762_  & \new_Sorter100|17763_ ;
  assign \new_Sorter100|17863_  = \new_Sorter100|17762_  | \new_Sorter100|17763_ ;
  assign \new_Sorter100|17864_  = \new_Sorter100|17764_  & \new_Sorter100|17765_ ;
  assign \new_Sorter100|17865_  = \new_Sorter100|17764_  | \new_Sorter100|17765_ ;
  assign \new_Sorter100|17866_  = \new_Sorter100|17766_  & \new_Sorter100|17767_ ;
  assign \new_Sorter100|17867_  = \new_Sorter100|17766_  | \new_Sorter100|17767_ ;
  assign \new_Sorter100|17868_  = \new_Sorter100|17768_  & \new_Sorter100|17769_ ;
  assign \new_Sorter100|17869_  = \new_Sorter100|17768_  | \new_Sorter100|17769_ ;
  assign \new_Sorter100|17870_  = \new_Sorter100|17770_  & \new_Sorter100|17771_ ;
  assign \new_Sorter100|17871_  = \new_Sorter100|17770_  | \new_Sorter100|17771_ ;
  assign \new_Sorter100|17872_  = \new_Sorter100|17772_  & \new_Sorter100|17773_ ;
  assign \new_Sorter100|17873_  = \new_Sorter100|17772_  | \new_Sorter100|17773_ ;
  assign \new_Sorter100|17874_  = \new_Sorter100|17774_  & \new_Sorter100|17775_ ;
  assign \new_Sorter100|17875_  = \new_Sorter100|17774_  | \new_Sorter100|17775_ ;
  assign \new_Sorter100|17876_  = \new_Sorter100|17776_  & \new_Sorter100|17777_ ;
  assign \new_Sorter100|17877_  = \new_Sorter100|17776_  | \new_Sorter100|17777_ ;
  assign \new_Sorter100|17878_  = \new_Sorter100|17778_  & \new_Sorter100|17779_ ;
  assign \new_Sorter100|17879_  = \new_Sorter100|17778_  | \new_Sorter100|17779_ ;
  assign \new_Sorter100|17880_  = \new_Sorter100|17780_  & \new_Sorter100|17781_ ;
  assign \new_Sorter100|17881_  = \new_Sorter100|17780_  | \new_Sorter100|17781_ ;
  assign \new_Sorter100|17882_  = \new_Sorter100|17782_  & \new_Sorter100|17783_ ;
  assign \new_Sorter100|17883_  = \new_Sorter100|17782_  | \new_Sorter100|17783_ ;
  assign \new_Sorter100|17884_  = \new_Sorter100|17784_  & \new_Sorter100|17785_ ;
  assign \new_Sorter100|17885_  = \new_Sorter100|17784_  | \new_Sorter100|17785_ ;
  assign \new_Sorter100|17886_  = \new_Sorter100|17786_  & \new_Sorter100|17787_ ;
  assign \new_Sorter100|17887_  = \new_Sorter100|17786_  | \new_Sorter100|17787_ ;
  assign \new_Sorter100|17888_  = \new_Sorter100|17788_  & \new_Sorter100|17789_ ;
  assign \new_Sorter100|17889_  = \new_Sorter100|17788_  | \new_Sorter100|17789_ ;
  assign \new_Sorter100|17890_  = \new_Sorter100|17790_  & \new_Sorter100|17791_ ;
  assign \new_Sorter100|17891_  = \new_Sorter100|17790_  | \new_Sorter100|17791_ ;
  assign \new_Sorter100|17892_  = \new_Sorter100|17792_  & \new_Sorter100|17793_ ;
  assign \new_Sorter100|17893_  = \new_Sorter100|17792_  | \new_Sorter100|17793_ ;
  assign \new_Sorter100|17894_  = \new_Sorter100|17794_  & \new_Sorter100|17795_ ;
  assign \new_Sorter100|17895_  = \new_Sorter100|17794_  | \new_Sorter100|17795_ ;
  assign \new_Sorter100|17896_  = \new_Sorter100|17796_  & \new_Sorter100|17797_ ;
  assign \new_Sorter100|17897_  = \new_Sorter100|17796_  | \new_Sorter100|17797_ ;
  assign \new_Sorter100|17898_  = \new_Sorter100|17798_  & \new_Sorter100|17799_ ;
  assign \new_Sorter100|17899_  = \new_Sorter100|17798_  | \new_Sorter100|17799_ ;
  assign \new_Sorter100|17900_  = \new_Sorter100|17800_ ;
  assign \new_Sorter100|17999_  = \new_Sorter100|17899_ ;
  assign \new_Sorter100|17901_  = \new_Sorter100|17801_  & \new_Sorter100|17802_ ;
  assign \new_Sorter100|17902_  = \new_Sorter100|17801_  | \new_Sorter100|17802_ ;
  assign \new_Sorter100|17903_  = \new_Sorter100|17803_  & \new_Sorter100|17804_ ;
  assign \new_Sorter100|17904_  = \new_Sorter100|17803_  | \new_Sorter100|17804_ ;
  assign \new_Sorter100|17905_  = \new_Sorter100|17805_  & \new_Sorter100|17806_ ;
  assign \new_Sorter100|17906_  = \new_Sorter100|17805_  | \new_Sorter100|17806_ ;
  assign \new_Sorter100|17907_  = \new_Sorter100|17807_  & \new_Sorter100|17808_ ;
  assign \new_Sorter100|17908_  = \new_Sorter100|17807_  | \new_Sorter100|17808_ ;
  assign \new_Sorter100|17909_  = \new_Sorter100|17809_  & \new_Sorter100|17810_ ;
  assign \new_Sorter100|17910_  = \new_Sorter100|17809_  | \new_Sorter100|17810_ ;
  assign \new_Sorter100|17911_  = \new_Sorter100|17811_  & \new_Sorter100|17812_ ;
  assign \new_Sorter100|17912_  = \new_Sorter100|17811_  | \new_Sorter100|17812_ ;
  assign \new_Sorter100|17913_  = \new_Sorter100|17813_  & \new_Sorter100|17814_ ;
  assign \new_Sorter100|17914_  = \new_Sorter100|17813_  | \new_Sorter100|17814_ ;
  assign \new_Sorter100|17915_  = \new_Sorter100|17815_  & \new_Sorter100|17816_ ;
  assign \new_Sorter100|17916_  = \new_Sorter100|17815_  | \new_Sorter100|17816_ ;
  assign \new_Sorter100|17917_  = \new_Sorter100|17817_  & \new_Sorter100|17818_ ;
  assign \new_Sorter100|17918_  = \new_Sorter100|17817_  | \new_Sorter100|17818_ ;
  assign \new_Sorter100|17919_  = \new_Sorter100|17819_  & \new_Sorter100|17820_ ;
  assign \new_Sorter100|17920_  = \new_Sorter100|17819_  | \new_Sorter100|17820_ ;
  assign \new_Sorter100|17921_  = \new_Sorter100|17821_  & \new_Sorter100|17822_ ;
  assign \new_Sorter100|17922_  = \new_Sorter100|17821_  | \new_Sorter100|17822_ ;
  assign \new_Sorter100|17923_  = \new_Sorter100|17823_  & \new_Sorter100|17824_ ;
  assign \new_Sorter100|17924_  = \new_Sorter100|17823_  | \new_Sorter100|17824_ ;
  assign \new_Sorter100|17925_  = \new_Sorter100|17825_  & \new_Sorter100|17826_ ;
  assign \new_Sorter100|17926_  = \new_Sorter100|17825_  | \new_Sorter100|17826_ ;
  assign \new_Sorter100|17927_  = \new_Sorter100|17827_  & \new_Sorter100|17828_ ;
  assign \new_Sorter100|17928_  = \new_Sorter100|17827_  | \new_Sorter100|17828_ ;
  assign \new_Sorter100|17929_  = \new_Sorter100|17829_  & \new_Sorter100|17830_ ;
  assign \new_Sorter100|17930_  = \new_Sorter100|17829_  | \new_Sorter100|17830_ ;
  assign \new_Sorter100|17931_  = \new_Sorter100|17831_  & \new_Sorter100|17832_ ;
  assign \new_Sorter100|17932_  = \new_Sorter100|17831_  | \new_Sorter100|17832_ ;
  assign \new_Sorter100|17933_  = \new_Sorter100|17833_  & \new_Sorter100|17834_ ;
  assign \new_Sorter100|17934_  = \new_Sorter100|17833_  | \new_Sorter100|17834_ ;
  assign \new_Sorter100|17935_  = \new_Sorter100|17835_  & \new_Sorter100|17836_ ;
  assign \new_Sorter100|17936_  = \new_Sorter100|17835_  | \new_Sorter100|17836_ ;
  assign \new_Sorter100|17937_  = \new_Sorter100|17837_  & \new_Sorter100|17838_ ;
  assign \new_Sorter100|17938_  = \new_Sorter100|17837_  | \new_Sorter100|17838_ ;
  assign \new_Sorter100|17939_  = \new_Sorter100|17839_  & \new_Sorter100|17840_ ;
  assign \new_Sorter100|17940_  = \new_Sorter100|17839_  | \new_Sorter100|17840_ ;
  assign \new_Sorter100|17941_  = \new_Sorter100|17841_  & \new_Sorter100|17842_ ;
  assign \new_Sorter100|17942_  = \new_Sorter100|17841_  | \new_Sorter100|17842_ ;
  assign \new_Sorter100|17943_  = \new_Sorter100|17843_  & \new_Sorter100|17844_ ;
  assign \new_Sorter100|17944_  = \new_Sorter100|17843_  | \new_Sorter100|17844_ ;
  assign \new_Sorter100|17945_  = \new_Sorter100|17845_  & \new_Sorter100|17846_ ;
  assign \new_Sorter100|17946_  = \new_Sorter100|17845_  | \new_Sorter100|17846_ ;
  assign \new_Sorter100|17947_  = \new_Sorter100|17847_  & \new_Sorter100|17848_ ;
  assign \new_Sorter100|17948_  = \new_Sorter100|17847_  | \new_Sorter100|17848_ ;
  assign \new_Sorter100|17949_  = \new_Sorter100|17849_  & \new_Sorter100|17850_ ;
  assign \new_Sorter100|17950_  = \new_Sorter100|17849_  | \new_Sorter100|17850_ ;
  assign \new_Sorter100|17951_  = \new_Sorter100|17851_  & \new_Sorter100|17852_ ;
  assign \new_Sorter100|17952_  = \new_Sorter100|17851_  | \new_Sorter100|17852_ ;
  assign \new_Sorter100|17953_  = \new_Sorter100|17853_  & \new_Sorter100|17854_ ;
  assign \new_Sorter100|17954_  = \new_Sorter100|17853_  | \new_Sorter100|17854_ ;
  assign \new_Sorter100|17955_  = \new_Sorter100|17855_  & \new_Sorter100|17856_ ;
  assign \new_Sorter100|17956_  = \new_Sorter100|17855_  | \new_Sorter100|17856_ ;
  assign \new_Sorter100|17957_  = \new_Sorter100|17857_  & \new_Sorter100|17858_ ;
  assign \new_Sorter100|17958_  = \new_Sorter100|17857_  | \new_Sorter100|17858_ ;
  assign \new_Sorter100|17959_  = \new_Sorter100|17859_  & \new_Sorter100|17860_ ;
  assign \new_Sorter100|17960_  = \new_Sorter100|17859_  | \new_Sorter100|17860_ ;
  assign \new_Sorter100|17961_  = \new_Sorter100|17861_  & \new_Sorter100|17862_ ;
  assign \new_Sorter100|17962_  = \new_Sorter100|17861_  | \new_Sorter100|17862_ ;
  assign \new_Sorter100|17963_  = \new_Sorter100|17863_  & \new_Sorter100|17864_ ;
  assign \new_Sorter100|17964_  = \new_Sorter100|17863_  | \new_Sorter100|17864_ ;
  assign \new_Sorter100|17965_  = \new_Sorter100|17865_  & \new_Sorter100|17866_ ;
  assign \new_Sorter100|17966_  = \new_Sorter100|17865_  | \new_Sorter100|17866_ ;
  assign \new_Sorter100|17967_  = \new_Sorter100|17867_  & \new_Sorter100|17868_ ;
  assign \new_Sorter100|17968_  = \new_Sorter100|17867_  | \new_Sorter100|17868_ ;
  assign \new_Sorter100|17969_  = \new_Sorter100|17869_  & \new_Sorter100|17870_ ;
  assign \new_Sorter100|17970_  = \new_Sorter100|17869_  | \new_Sorter100|17870_ ;
  assign \new_Sorter100|17971_  = \new_Sorter100|17871_  & \new_Sorter100|17872_ ;
  assign \new_Sorter100|17972_  = \new_Sorter100|17871_  | \new_Sorter100|17872_ ;
  assign \new_Sorter100|17973_  = \new_Sorter100|17873_  & \new_Sorter100|17874_ ;
  assign \new_Sorter100|17974_  = \new_Sorter100|17873_  | \new_Sorter100|17874_ ;
  assign \new_Sorter100|17975_  = \new_Sorter100|17875_  & \new_Sorter100|17876_ ;
  assign \new_Sorter100|17976_  = \new_Sorter100|17875_  | \new_Sorter100|17876_ ;
  assign \new_Sorter100|17977_  = \new_Sorter100|17877_  & \new_Sorter100|17878_ ;
  assign \new_Sorter100|17978_  = \new_Sorter100|17877_  | \new_Sorter100|17878_ ;
  assign \new_Sorter100|17979_  = \new_Sorter100|17879_  & \new_Sorter100|17880_ ;
  assign \new_Sorter100|17980_  = \new_Sorter100|17879_  | \new_Sorter100|17880_ ;
  assign \new_Sorter100|17981_  = \new_Sorter100|17881_  & \new_Sorter100|17882_ ;
  assign \new_Sorter100|17982_  = \new_Sorter100|17881_  | \new_Sorter100|17882_ ;
  assign \new_Sorter100|17983_  = \new_Sorter100|17883_  & \new_Sorter100|17884_ ;
  assign \new_Sorter100|17984_  = \new_Sorter100|17883_  | \new_Sorter100|17884_ ;
  assign \new_Sorter100|17985_  = \new_Sorter100|17885_  & \new_Sorter100|17886_ ;
  assign \new_Sorter100|17986_  = \new_Sorter100|17885_  | \new_Sorter100|17886_ ;
  assign \new_Sorter100|17987_  = \new_Sorter100|17887_  & \new_Sorter100|17888_ ;
  assign \new_Sorter100|17988_  = \new_Sorter100|17887_  | \new_Sorter100|17888_ ;
  assign \new_Sorter100|17989_  = \new_Sorter100|17889_  & \new_Sorter100|17890_ ;
  assign \new_Sorter100|17990_  = \new_Sorter100|17889_  | \new_Sorter100|17890_ ;
  assign \new_Sorter100|17991_  = \new_Sorter100|17891_  & \new_Sorter100|17892_ ;
  assign \new_Sorter100|17992_  = \new_Sorter100|17891_  | \new_Sorter100|17892_ ;
  assign \new_Sorter100|17993_  = \new_Sorter100|17893_  & \new_Sorter100|17894_ ;
  assign \new_Sorter100|17994_  = \new_Sorter100|17893_  | \new_Sorter100|17894_ ;
  assign \new_Sorter100|17995_  = \new_Sorter100|17895_  & \new_Sorter100|17896_ ;
  assign \new_Sorter100|17996_  = \new_Sorter100|17895_  | \new_Sorter100|17896_ ;
  assign \new_Sorter100|17997_  = \new_Sorter100|17897_  & \new_Sorter100|17898_ ;
  assign \new_Sorter100|17998_  = \new_Sorter100|17897_  | \new_Sorter100|17898_ ;
  assign \new_Sorter100|18000_  = \new_Sorter100|17900_  & \new_Sorter100|17901_ ;
  assign \new_Sorter100|18001_  = \new_Sorter100|17900_  | \new_Sorter100|17901_ ;
  assign \new_Sorter100|18002_  = \new_Sorter100|17902_  & \new_Sorter100|17903_ ;
  assign \new_Sorter100|18003_  = \new_Sorter100|17902_  | \new_Sorter100|17903_ ;
  assign \new_Sorter100|18004_  = \new_Sorter100|17904_  & \new_Sorter100|17905_ ;
  assign \new_Sorter100|18005_  = \new_Sorter100|17904_  | \new_Sorter100|17905_ ;
  assign \new_Sorter100|18006_  = \new_Sorter100|17906_  & \new_Sorter100|17907_ ;
  assign \new_Sorter100|18007_  = \new_Sorter100|17906_  | \new_Sorter100|17907_ ;
  assign \new_Sorter100|18008_  = \new_Sorter100|17908_  & \new_Sorter100|17909_ ;
  assign \new_Sorter100|18009_  = \new_Sorter100|17908_  | \new_Sorter100|17909_ ;
  assign \new_Sorter100|18010_  = \new_Sorter100|17910_  & \new_Sorter100|17911_ ;
  assign \new_Sorter100|18011_  = \new_Sorter100|17910_  | \new_Sorter100|17911_ ;
  assign \new_Sorter100|18012_  = \new_Sorter100|17912_  & \new_Sorter100|17913_ ;
  assign \new_Sorter100|18013_  = \new_Sorter100|17912_  | \new_Sorter100|17913_ ;
  assign \new_Sorter100|18014_  = \new_Sorter100|17914_  & \new_Sorter100|17915_ ;
  assign \new_Sorter100|18015_  = \new_Sorter100|17914_  | \new_Sorter100|17915_ ;
  assign \new_Sorter100|18016_  = \new_Sorter100|17916_  & \new_Sorter100|17917_ ;
  assign \new_Sorter100|18017_  = \new_Sorter100|17916_  | \new_Sorter100|17917_ ;
  assign \new_Sorter100|18018_  = \new_Sorter100|17918_  & \new_Sorter100|17919_ ;
  assign \new_Sorter100|18019_  = \new_Sorter100|17918_  | \new_Sorter100|17919_ ;
  assign \new_Sorter100|18020_  = \new_Sorter100|17920_  & \new_Sorter100|17921_ ;
  assign \new_Sorter100|18021_  = \new_Sorter100|17920_  | \new_Sorter100|17921_ ;
  assign \new_Sorter100|18022_  = \new_Sorter100|17922_  & \new_Sorter100|17923_ ;
  assign \new_Sorter100|18023_  = \new_Sorter100|17922_  | \new_Sorter100|17923_ ;
  assign \new_Sorter100|18024_  = \new_Sorter100|17924_  & \new_Sorter100|17925_ ;
  assign \new_Sorter100|18025_  = \new_Sorter100|17924_  | \new_Sorter100|17925_ ;
  assign \new_Sorter100|18026_  = \new_Sorter100|17926_  & \new_Sorter100|17927_ ;
  assign \new_Sorter100|18027_  = \new_Sorter100|17926_  | \new_Sorter100|17927_ ;
  assign \new_Sorter100|18028_  = \new_Sorter100|17928_  & \new_Sorter100|17929_ ;
  assign \new_Sorter100|18029_  = \new_Sorter100|17928_  | \new_Sorter100|17929_ ;
  assign \new_Sorter100|18030_  = \new_Sorter100|17930_  & \new_Sorter100|17931_ ;
  assign \new_Sorter100|18031_  = \new_Sorter100|17930_  | \new_Sorter100|17931_ ;
  assign \new_Sorter100|18032_  = \new_Sorter100|17932_  & \new_Sorter100|17933_ ;
  assign \new_Sorter100|18033_  = \new_Sorter100|17932_  | \new_Sorter100|17933_ ;
  assign \new_Sorter100|18034_  = \new_Sorter100|17934_  & \new_Sorter100|17935_ ;
  assign \new_Sorter100|18035_  = \new_Sorter100|17934_  | \new_Sorter100|17935_ ;
  assign \new_Sorter100|18036_  = \new_Sorter100|17936_  & \new_Sorter100|17937_ ;
  assign \new_Sorter100|18037_  = \new_Sorter100|17936_  | \new_Sorter100|17937_ ;
  assign \new_Sorter100|18038_  = \new_Sorter100|17938_  & \new_Sorter100|17939_ ;
  assign \new_Sorter100|18039_  = \new_Sorter100|17938_  | \new_Sorter100|17939_ ;
  assign \new_Sorter100|18040_  = \new_Sorter100|17940_  & \new_Sorter100|17941_ ;
  assign \new_Sorter100|18041_  = \new_Sorter100|17940_  | \new_Sorter100|17941_ ;
  assign \new_Sorter100|18042_  = \new_Sorter100|17942_  & \new_Sorter100|17943_ ;
  assign \new_Sorter100|18043_  = \new_Sorter100|17942_  | \new_Sorter100|17943_ ;
  assign \new_Sorter100|18044_  = \new_Sorter100|17944_  & \new_Sorter100|17945_ ;
  assign \new_Sorter100|18045_  = \new_Sorter100|17944_  | \new_Sorter100|17945_ ;
  assign \new_Sorter100|18046_  = \new_Sorter100|17946_  & \new_Sorter100|17947_ ;
  assign \new_Sorter100|18047_  = \new_Sorter100|17946_  | \new_Sorter100|17947_ ;
  assign \new_Sorter100|18048_  = \new_Sorter100|17948_  & \new_Sorter100|17949_ ;
  assign \new_Sorter100|18049_  = \new_Sorter100|17948_  | \new_Sorter100|17949_ ;
  assign \new_Sorter100|18050_  = \new_Sorter100|17950_  & \new_Sorter100|17951_ ;
  assign \new_Sorter100|18051_  = \new_Sorter100|17950_  | \new_Sorter100|17951_ ;
  assign \new_Sorter100|18052_  = \new_Sorter100|17952_  & \new_Sorter100|17953_ ;
  assign \new_Sorter100|18053_  = \new_Sorter100|17952_  | \new_Sorter100|17953_ ;
  assign \new_Sorter100|18054_  = \new_Sorter100|17954_  & \new_Sorter100|17955_ ;
  assign \new_Sorter100|18055_  = \new_Sorter100|17954_  | \new_Sorter100|17955_ ;
  assign \new_Sorter100|18056_  = \new_Sorter100|17956_  & \new_Sorter100|17957_ ;
  assign \new_Sorter100|18057_  = \new_Sorter100|17956_  | \new_Sorter100|17957_ ;
  assign \new_Sorter100|18058_  = \new_Sorter100|17958_  & \new_Sorter100|17959_ ;
  assign \new_Sorter100|18059_  = \new_Sorter100|17958_  | \new_Sorter100|17959_ ;
  assign \new_Sorter100|18060_  = \new_Sorter100|17960_  & \new_Sorter100|17961_ ;
  assign \new_Sorter100|18061_  = \new_Sorter100|17960_  | \new_Sorter100|17961_ ;
  assign \new_Sorter100|18062_  = \new_Sorter100|17962_  & \new_Sorter100|17963_ ;
  assign \new_Sorter100|18063_  = \new_Sorter100|17962_  | \new_Sorter100|17963_ ;
  assign \new_Sorter100|18064_  = \new_Sorter100|17964_  & \new_Sorter100|17965_ ;
  assign \new_Sorter100|18065_  = \new_Sorter100|17964_  | \new_Sorter100|17965_ ;
  assign \new_Sorter100|18066_  = \new_Sorter100|17966_  & \new_Sorter100|17967_ ;
  assign \new_Sorter100|18067_  = \new_Sorter100|17966_  | \new_Sorter100|17967_ ;
  assign \new_Sorter100|18068_  = \new_Sorter100|17968_  & \new_Sorter100|17969_ ;
  assign \new_Sorter100|18069_  = \new_Sorter100|17968_  | \new_Sorter100|17969_ ;
  assign \new_Sorter100|18070_  = \new_Sorter100|17970_  & \new_Sorter100|17971_ ;
  assign \new_Sorter100|18071_  = \new_Sorter100|17970_  | \new_Sorter100|17971_ ;
  assign \new_Sorter100|18072_  = \new_Sorter100|17972_  & \new_Sorter100|17973_ ;
  assign \new_Sorter100|18073_  = \new_Sorter100|17972_  | \new_Sorter100|17973_ ;
  assign \new_Sorter100|18074_  = \new_Sorter100|17974_  & \new_Sorter100|17975_ ;
  assign \new_Sorter100|18075_  = \new_Sorter100|17974_  | \new_Sorter100|17975_ ;
  assign \new_Sorter100|18076_  = \new_Sorter100|17976_  & \new_Sorter100|17977_ ;
  assign \new_Sorter100|18077_  = \new_Sorter100|17976_  | \new_Sorter100|17977_ ;
  assign \new_Sorter100|18078_  = \new_Sorter100|17978_  & \new_Sorter100|17979_ ;
  assign \new_Sorter100|18079_  = \new_Sorter100|17978_  | \new_Sorter100|17979_ ;
  assign \new_Sorter100|18080_  = \new_Sorter100|17980_  & \new_Sorter100|17981_ ;
  assign \new_Sorter100|18081_  = \new_Sorter100|17980_  | \new_Sorter100|17981_ ;
  assign \new_Sorter100|18082_  = \new_Sorter100|17982_  & \new_Sorter100|17983_ ;
  assign \new_Sorter100|18083_  = \new_Sorter100|17982_  | \new_Sorter100|17983_ ;
  assign \new_Sorter100|18084_  = \new_Sorter100|17984_  & \new_Sorter100|17985_ ;
  assign \new_Sorter100|18085_  = \new_Sorter100|17984_  | \new_Sorter100|17985_ ;
  assign \new_Sorter100|18086_  = \new_Sorter100|17986_  & \new_Sorter100|17987_ ;
  assign \new_Sorter100|18087_  = \new_Sorter100|17986_  | \new_Sorter100|17987_ ;
  assign \new_Sorter100|18088_  = \new_Sorter100|17988_  & \new_Sorter100|17989_ ;
  assign \new_Sorter100|18089_  = \new_Sorter100|17988_  | \new_Sorter100|17989_ ;
  assign \new_Sorter100|18090_  = \new_Sorter100|17990_  & \new_Sorter100|17991_ ;
  assign \new_Sorter100|18091_  = \new_Sorter100|17990_  | \new_Sorter100|17991_ ;
  assign \new_Sorter100|18092_  = \new_Sorter100|17992_  & \new_Sorter100|17993_ ;
  assign \new_Sorter100|18093_  = \new_Sorter100|17992_  | \new_Sorter100|17993_ ;
  assign \new_Sorter100|18094_  = \new_Sorter100|17994_  & \new_Sorter100|17995_ ;
  assign \new_Sorter100|18095_  = \new_Sorter100|17994_  | \new_Sorter100|17995_ ;
  assign \new_Sorter100|18096_  = \new_Sorter100|17996_  & \new_Sorter100|17997_ ;
  assign \new_Sorter100|18097_  = \new_Sorter100|17996_  | \new_Sorter100|17997_ ;
  assign \new_Sorter100|18098_  = \new_Sorter100|17998_  & \new_Sorter100|17999_ ;
  assign \new_Sorter100|18099_  = \new_Sorter100|17998_  | \new_Sorter100|17999_ ;
  assign \new_Sorter100|18100_  = \new_Sorter100|18000_ ;
  assign \new_Sorter100|18199_  = \new_Sorter100|18099_ ;
  assign \new_Sorter100|18101_  = \new_Sorter100|18001_  & \new_Sorter100|18002_ ;
  assign \new_Sorter100|18102_  = \new_Sorter100|18001_  | \new_Sorter100|18002_ ;
  assign \new_Sorter100|18103_  = \new_Sorter100|18003_  & \new_Sorter100|18004_ ;
  assign \new_Sorter100|18104_  = \new_Sorter100|18003_  | \new_Sorter100|18004_ ;
  assign \new_Sorter100|18105_  = \new_Sorter100|18005_  & \new_Sorter100|18006_ ;
  assign \new_Sorter100|18106_  = \new_Sorter100|18005_  | \new_Sorter100|18006_ ;
  assign \new_Sorter100|18107_  = \new_Sorter100|18007_  & \new_Sorter100|18008_ ;
  assign \new_Sorter100|18108_  = \new_Sorter100|18007_  | \new_Sorter100|18008_ ;
  assign \new_Sorter100|18109_  = \new_Sorter100|18009_  & \new_Sorter100|18010_ ;
  assign \new_Sorter100|18110_  = \new_Sorter100|18009_  | \new_Sorter100|18010_ ;
  assign \new_Sorter100|18111_  = \new_Sorter100|18011_  & \new_Sorter100|18012_ ;
  assign \new_Sorter100|18112_  = \new_Sorter100|18011_  | \new_Sorter100|18012_ ;
  assign \new_Sorter100|18113_  = \new_Sorter100|18013_  & \new_Sorter100|18014_ ;
  assign \new_Sorter100|18114_  = \new_Sorter100|18013_  | \new_Sorter100|18014_ ;
  assign \new_Sorter100|18115_  = \new_Sorter100|18015_  & \new_Sorter100|18016_ ;
  assign \new_Sorter100|18116_  = \new_Sorter100|18015_  | \new_Sorter100|18016_ ;
  assign \new_Sorter100|18117_  = \new_Sorter100|18017_  & \new_Sorter100|18018_ ;
  assign \new_Sorter100|18118_  = \new_Sorter100|18017_  | \new_Sorter100|18018_ ;
  assign \new_Sorter100|18119_  = \new_Sorter100|18019_  & \new_Sorter100|18020_ ;
  assign \new_Sorter100|18120_  = \new_Sorter100|18019_  | \new_Sorter100|18020_ ;
  assign \new_Sorter100|18121_  = \new_Sorter100|18021_  & \new_Sorter100|18022_ ;
  assign \new_Sorter100|18122_  = \new_Sorter100|18021_  | \new_Sorter100|18022_ ;
  assign \new_Sorter100|18123_  = \new_Sorter100|18023_  & \new_Sorter100|18024_ ;
  assign \new_Sorter100|18124_  = \new_Sorter100|18023_  | \new_Sorter100|18024_ ;
  assign \new_Sorter100|18125_  = \new_Sorter100|18025_  & \new_Sorter100|18026_ ;
  assign \new_Sorter100|18126_  = \new_Sorter100|18025_  | \new_Sorter100|18026_ ;
  assign \new_Sorter100|18127_  = \new_Sorter100|18027_  & \new_Sorter100|18028_ ;
  assign \new_Sorter100|18128_  = \new_Sorter100|18027_  | \new_Sorter100|18028_ ;
  assign \new_Sorter100|18129_  = \new_Sorter100|18029_  & \new_Sorter100|18030_ ;
  assign \new_Sorter100|18130_  = \new_Sorter100|18029_  | \new_Sorter100|18030_ ;
  assign \new_Sorter100|18131_  = \new_Sorter100|18031_  & \new_Sorter100|18032_ ;
  assign \new_Sorter100|18132_  = \new_Sorter100|18031_  | \new_Sorter100|18032_ ;
  assign \new_Sorter100|18133_  = \new_Sorter100|18033_  & \new_Sorter100|18034_ ;
  assign \new_Sorter100|18134_  = \new_Sorter100|18033_  | \new_Sorter100|18034_ ;
  assign \new_Sorter100|18135_  = \new_Sorter100|18035_  & \new_Sorter100|18036_ ;
  assign \new_Sorter100|18136_  = \new_Sorter100|18035_  | \new_Sorter100|18036_ ;
  assign \new_Sorter100|18137_  = \new_Sorter100|18037_  & \new_Sorter100|18038_ ;
  assign \new_Sorter100|18138_  = \new_Sorter100|18037_  | \new_Sorter100|18038_ ;
  assign \new_Sorter100|18139_  = \new_Sorter100|18039_  & \new_Sorter100|18040_ ;
  assign \new_Sorter100|18140_  = \new_Sorter100|18039_  | \new_Sorter100|18040_ ;
  assign \new_Sorter100|18141_  = \new_Sorter100|18041_  & \new_Sorter100|18042_ ;
  assign \new_Sorter100|18142_  = \new_Sorter100|18041_  | \new_Sorter100|18042_ ;
  assign \new_Sorter100|18143_  = \new_Sorter100|18043_  & \new_Sorter100|18044_ ;
  assign \new_Sorter100|18144_  = \new_Sorter100|18043_  | \new_Sorter100|18044_ ;
  assign \new_Sorter100|18145_  = \new_Sorter100|18045_  & \new_Sorter100|18046_ ;
  assign \new_Sorter100|18146_  = \new_Sorter100|18045_  | \new_Sorter100|18046_ ;
  assign \new_Sorter100|18147_  = \new_Sorter100|18047_  & \new_Sorter100|18048_ ;
  assign \new_Sorter100|18148_  = \new_Sorter100|18047_  | \new_Sorter100|18048_ ;
  assign \new_Sorter100|18149_  = \new_Sorter100|18049_  & \new_Sorter100|18050_ ;
  assign \new_Sorter100|18150_  = \new_Sorter100|18049_  | \new_Sorter100|18050_ ;
  assign \new_Sorter100|18151_  = \new_Sorter100|18051_  & \new_Sorter100|18052_ ;
  assign \new_Sorter100|18152_  = \new_Sorter100|18051_  | \new_Sorter100|18052_ ;
  assign \new_Sorter100|18153_  = \new_Sorter100|18053_  & \new_Sorter100|18054_ ;
  assign \new_Sorter100|18154_  = \new_Sorter100|18053_  | \new_Sorter100|18054_ ;
  assign \new_Sorter100|18155_  = \new_Sorter100|18055_  & \new_Sorter100|18056_ ;
  assign \new_Sorter100|18156_  = \new_Sorter100|18055_  | \new_Sorter100|18056_ ;
  assign \new_Sorter100|18157_  = \new_Sorter100|18057_  & \new_Sorter100|18058_ ;
  assign \new_Sorter100|18158_  = \new_Sorter100|18057_  | \new_Sorter100|18058_ ;
  assign \new_Sorter100|18159_  = \new_Sorter100|18059_  & \new_Sorter100|18060_ ;
  assign \new_Sorter100|18160_  = \new_Sorter100|18059_  | \new_Sorter100|18060_ ;
  assign \new_Sorter100|18161_  = \new_Sorter100|18061_  & \new_Sorter100|18062_ ;
  assign \new_Sorter100|18162_  = \new_Sorter100|18061_  | \new_Sorter100|18062_ ;
  assign \new_Sorter100|18163_  = \new_Sorter100|18063_  & \new_Sorter100|18064_ ;
  assign \new_Sorter100|18164_  = \new_Sorter100|18063_  | \new_Sorter100|18064_ ;
  assign \new_Sorter100|18165_  = \new_Sorter100|18065_  & \new_Sorter100|18066_ ;
  assign \new_Sorter100|18166_  = \new_Sorter100|18065_  | \new_Sorter100|18066_ ;
  assign \new_Sorter100|18167_  = \new_Sorter100|18067_  & \new_Sorter100|18068_ ;
  assign \new_Sorter100|18168_  = \new_Sorter100|18067_  | \new_Sorter100|18068_ ;
  assign \new_Sorter100|18169_  = \new_Sorter100|18069_  & \new_Sorter100|18070_ ;
  assign \new_Sorter100|18170_  = \new_Sorter100|18069_  | \new_Sorter100|18070_ ;
  assign \new_Sorter100|18171_  = \new_Sorter100|18071_  & \new_Sorter100|18072_ ;
  assign \new_Sorter100|18172_  = \new_Sorter100|18071_  | \new_Sorter100|18072_ ;
  assign \new_Sorter100|18173_  = \new_Sorter100|18073_  & \new_Sorter100|18074_ ;
  assign \new_Sorter100|18174_  = \new_Sorter100|18073_  | \new_Sorter100|18074_ ;
  assign \new_Sorter100|18175_  = \new_Sorter100|18075_  & \new_Sorter100|18076_ ;
  assign \new_Sorter100|18176_  = \new_Sorter100|18075_  | \new_Sorter100|18076_ ;
  assign \new_Sorter100|18177_  = \new_Sorter100|18077_  & \new_Sorter100|18078_ ;
  assign \new_Sorter100|18178_  = \new_Sorter100|18077_  | \new_Sorter100|18078_ ;
  assign \new_Sorter100|18179_  = \new_Sorter100|18079_  & \new_Sorter100|18080_ ;
  assign \new_Sorter100|18180_  = \new_Sorter100|18079_  | \new_Sorter100|18080_ ;
  assign \new_Sorter100|18181_  = \new_Sorter100|18081_  & \new_Sorter100|18082_ ;
  assign \new_Sorter100|18182_  = \new_Sorter100|18081_  | \new_Sorter100|18082_ ;
  assign \new_Sorter100|18183_  = \new_Sorter100|18083_  & \new_Sorter100|18084_ ;
  assign \new_Sorter100|18184_  = \new_Sorter100|18083_  | \new_Sorter100|18084_ ;
  assign \new_Sorter100|18185_  = \new_Sorter100|18085_  & \new_Sorter100|18086_ ;
  assign \new_Sorter100|18186_  = \new_Sorter100|18085_  | \new_Sorter100|18086_ ;
  assign \new_Sorter100|18187_  = \new_Sorter100|18087_  & \new_Sorter100|18088_ ;
  assign \new_Sorter100|18188_  = \new_Sorter100|18087_  | \new_Sorter100|18088_ ;
  assign \new_Sorter100|18189_  = \new_Sorter100|18089_  & \new_Sorter100|18090_ ;
  assign \new_Sorter100|18190_  = \new_Sorter100|18089_  | \new_Sorter100|18090_ ;
  assign \new_Sorter100|18191_  = \new_Sorter100|18091_  & \new_Sorter100|18092_ ;
  assign \new_Sorter100|18192_  = \new_Sorter100|18091_  | \new_Sorter100|18092_ ;
  assign \new_Sorter100|18193_  = \new_Sorter100|18093_  & \new_Sorter100|18094_ ;
  assign \new_Sorter100|18194_  = \new_Sorter100|18093_  | \new_Sorter100|18094_ ;
  assign \new_Sorter100|18195_  = \new_Sorter100|18095_  & \new_Sorter100|18096_ ;
  assign \new_Sorter100|18196_  = \new_Sorter100|18095_  | \new_Sorter100|18096_ ;
  assign \new_Sorter100|18197_  = \new_Sorter100|18097_  & \new_Sorter100|18098_ ;
  assign \new_Sorter100|18198_  = \new_Sorter100|18097_  | \new_Sorter100|18098_ ;
  assign \new_Sorter100|18200_  = \new_Sorter100|18100_  & \new_Sorter100|18101_ ;
  assign \new_Sorter100|18201_  = \new_Sorter100|18100_  | \new_Sorter100|18101_ ;
  assign \new_Sorter100|18202_  = \new_Sorter100|18102_  & \new_Sorter100|18103_ ;
  assign \new_Sorter100|18203_  = \new_Sorter100|18102_  | \new_Sorter100|18103_ ;
  assign \new_Sorter100|18204_  = \new_Sorter100|18104_  & \new_Sorter100|18105_ ;
  assign \new_Sorter100|18205_  = \new_Sorter100|18104_  | \new_Sorter100|18105_ ;
  assign \new_Sorter100|18206_  = \new_Sorter100|18106_  & \new_Sorter100|18107_ ;
  assign \new_Sorter100|18207_  = \new_Sorter100|18106_  | \new_Sorter100|18107_ ;
  assign \new_Sorter100|18208_  = \new_Sorter100|18108_  & \new_Sorter100|18109_ ;
  assign \new_Sorter100|18209_  = \new_Sorter100|18108_  | \new_Sorter100|18109_ ;
  assign \new_Sorter100|18210_  = \new_Sorter100|18110_  & \new_Sorter100|18111_ ;
  assign \new_Sorter100|18211_  = \new_Sorter100|18110_  | \new_Sorter100|18111_ ;
  assign \new_Sorter100|18212_  = \new_Sorter100|18112_  & \new_Sorter100|18113_ ;
  assign \new_Sorter100|18213_  = \new_Sorter100|18112_  | \new_Sorter100|18113_ ;
  assign \new_Sorter100|18214_  = \new_Sorter100|18114_  & \new_Sorter100|18115_ ;
  assign \new_Sorter100|18215_  = \new_Sorter100|18114_  | \new_Sorter100|18115_ ;
  assign \new_Sorter100|18216_  = \new_Sorter100|18116_  & \new_Sorter100|18117_ ;
  assign \new_Sorter100|18217_  = \new_Sorter100|18116_  | \new_Sorter100|18117_ ;
  assign \new_Sorter100|18218_  = \new_Sorter100|18118_  & \new_Sorter100|18119_ ;
  assign \new_Sorter100|18219_  = \new_Sorter100|18118_  | \new_Sorter100|18119_ ;
  assign \new_Sorter100|18220_  = \new_Sorter100|18120_  & \new_Sorter100|18121_ ;
  assign \new_Sorter100|18221_  = \new_Sorter100|18120_  | \new_Sorter100|18121_ ;
  assign \new_Sorter100|18222_  = \new_Sorter100|18122_  & \new_Sorter100|18123_ ;
  assign \new_Sorter100|18223_  = \new_Sorter100|18122_  | \new_Sorter100|18123_ ;
  assign \new_Sorter100|18224_  = \new_Sorter100|18124_  & \new_Sorter100|18125_ ;
  assign \new_Sorter100|18225_  = \new_Sorter100|18124_  | \new_Sorter100|18125_ ;
  assign \new_Sorter100|18226_  = \new_Sorter100|18126_  & \new_Sorter100|18127_ ;
  assign \new_Sorter100|18227_  = \new_Sorter100|18126_  | \new_Sorter100|18127_ ;
  assign \new_Sorter100|18228_  = \new_Sorter100|18128_  & \new_Sorter100|18129_ ;
  assign \new_Sorter100|18229_  = \new_Sorter100|18128_  | \new_Sorter100|18129_ ;
  assign \new_Sorter100|18230_  = \new_Sorter100|18130_  & \new_Sorter100|18131_ ;
  assign \new_Sorter100|18231_  = \new_Sorter100|18130_  | \new_Sorter100|18131_ ;
  assign \new_Sorter100|18232_  = \new_Sorter100|18132_  & \new_Sorter100|18133_ ;
  assign \new_Sorter100|18233_  = \new_Sorter100|18132_  | \new_Sorter100|18133_ ;
  assign \new_Sorter100|18234_  = \new_Sorter100|18134_  & \new_Sorter100|18135_ ;
  assign \new_Sorter100|18235_  = \new_Sorter100|18134_  | \new_Sorter100|18135_ ;
  assign \new_Sorter100|18236_  = \new_Sorter100|18136_  & \new_Sorter100|18137_ ;
  assign \new_Sorter100|18237_  = \new_Sorter100|18136_  | \new_Sorter100|18137_ ;
  assign \new_Sorter100|18238_  = \new_Sorter100|18138_  & \new_Sorter100|18139_ ;
  assign \new_Sorter100|18239_  = \new_Sorter100|18138_  | \new_Sorter100|18139_ ;
  assign \new_Sorter100|18240_  = \new_Sorter100|18140_  & \new_Sorter100|18141_ ;
  assign \new_Sorter100|18241_  = \new_Sorter100|18140_  | \new_Sorter100|18141_ ;
  assign \new_Sorter100|18242_  = \new_Sorter100|18142_  & \new_Sorter100|18143_ ;
  assign \new_Sorter100|18243_  = \new_Sorter100|18142_  | \new_Sorter100|18143_ ;
  assign \new_Sorter100|18244_  = \new_Sorter100|18144_  & \new_Sorter100|18145_ ;
  assign \new_Sorter100|18245_  = \new_Sorter100|18144_  | \new_Sorter100|18145_ ;
  assign \new_Sorter100|18246_  = \new_Sorter100|18146_  & \new_Sorter100|18147_ ;
  assign \new_Sorter100|18247_  = \new_Sorter100|18146_  | \new_Sorter100|18147_ ;
  assign \new_Sorter100|18248_  = \new_Sorter100|18148_  & \new_Sorter100|18149_ ;
  assign \new_Sorter100|18249_  = \new_Sorter100|18148_  | \new_Sorter100|18149_ ;
  assign \new_Sorter100|18250_  = \new_Sorter100|18150_  & \new_Sorter100|18151_ ;
  assign \new_Sorter100|18251_  = \new_Sorter100|18150_  | \new_Sorter100|18151_ ;
  assign \new_Sorter100|18252_  = \new_Sorter100|18152_  & \new_Sorter100|18153_ ;
  assign \new_Sorter100|18253_  = \new_Sorter100|18152_  | \new_Sorter100|18153_ ;
  assign \new_Sorter100|18254_  = \new_Sorter100|18154_  & \new_Sorter100|18155_ ;
  assign \new_Sorter100|18255_  = \new_Sorter100|18154_  | \new_Sorter100|18155_ ;
  assign \new_Sorter100|18256_  = \new_Sorter100|18156_  & \new_Sorter100|18157_ ;
  assign \new_Sorter100|18257_  = \new_Sorter100|18156_  | \new_Sorter100|18157_ ;
  assign \new_Sorter100|18258_  = \new_Sorter100|18158_  & \new_Sorter100|18159_ ;
  assign \new_Sorter100|18259_  = \new_Sorter100|18158_  | \new_Sorter100|18159_ ;
  assign \new_Sorter100|18260_  = \new_Sorter100|18160_  & \new_Sorter100|18161_ ;
  assign \new_Sorter100|18261_  = \new_Sorter100|18160_  | \new_Sorter100|18161_ ;
  assign \new_Sorter100|18262_  = \new_Sorter100|18162_  & \new_Sorter100|18163_ ;
  assign \new_Sorter100|18263_  = \new_Sorter100|18162_  | \new_Sorter100|18163_ ;
  assign \new_Sorter100|18264_  = \new_Sorter100|18164_  & \new_Sorter100|18165_ ;
  assign \new_Sorter100|18265_  = \new_Sorter100|18164_  | \new_Sorter100|18165_ ;
  assign \new_Sorter100|18266_  = \new_Sorter100|18166_  & \new_Sorter100|18167_ ;
  assign \new_Sorter100|18267_  = \new_Sorter100|18166_  | \new_Sorter100|18167_ ;
  assign \new_Sorter100|18268_  = \new_Sorter100|18168_  & \new_Sorter100|18169_ ;
  assign \new_Sorter100|18269_  = \new_Sorter100|18168_  | \new_Sorter100|18169_ ;
  assign \new_Sorter100|18270_  = \new_Sorter100|18170_  & \new_Sorter100|18171_ ;
  assign \new_Sorter100|18271_  = \new_Sorter100|18170_  | \new_Sorter100|18171_ ;
  assign \new_Sorter100|18272_  = \new_Sorter100|18172_  & \new_Sorter100|18173_ ;
  assign \new_Sorter100|18273_  = \new_Sorter100|18172_  | \new_Sorter100|18173_ ;
  assign \new_Sorter100|18274_  = \new_Sorter100|18174_  & \new_Sorter100|18175_ ;
  assign \new_Sorter100|18275_  = \new_Sorter100|18174_  | \new_Sorter100|18175_ ;
  assign \new_Sorter100|18276_  = \new_Sorter100|18176_  & \new_Sorter100|18177_ ;
  assign \new_Sorter100|18277_  = \new_Sorter100|18176_  | \new_Sorter100|18177_ ;
  assign \new_Sorter100|18278_  = \new_Sorter100|18178_  & \new_Sorter100|18179_ ;
  assign \new_Sorter100|18279_  = \new_Sorter100|18178_  | \new_Sorter100|18179_ ;
  assign \new_Sorter100|18280_  = \new_Sorter100|18180_  & \new_Sorter100|18181_ ;
  assign \new_Sorter100|18281_  = \new_Sorter100|18180_  | \new_Sorter100|18181_ ;
  assign \new_Sorter100|18282_  = \new_Sorter100|18182_  & \new_Sorter100|18183_ ;
  assign \new_Sorter100|18283_  = \new_Sorter100|18182_  | \new_Sorter100|18183_ ;
  assign \new_Sorter100|18284_  = \new_Sorter100|18184_  & \new_Sorter100|18185_ ;
  assign \new_Sorter100|18285_  = \new_Sorter100|18184_  | \new_Sorter100|18185_ ;
  assign \new_Sorter100|18286_  = \new_Sorter100|18186_  & \new_Sorter100|18187_ ;
  assign \new_Sorter100|18287_  = \new_Sorter100|18186_  | \new_Sorter100|18187_ ;
  assign \new_Sorter100|18288_  = \new_Sorter100|18188_  & \new_Sorter100|18189_ ;
  assign \new_Sorter100|18289_  = \new_Sorter100|18188_  | \new_Sorter100|18189_ ;
  assign \new_Sorter100|18290_  = \new_Sorter100|18190_  & \new_Sorter100|18191_ ;
  assign \new_Sorter100|18291_  = \new_Sorter100|18190_  | \new_Sorter100|18191_ ;
  assign \new_Sorter100|18292_  = \new_Sorter100|18192_  & \new_Sorter100|18193_ ;
  assign \new_Sorter100|18293_  = \new_Sorter100|18192_  | \new_Sorter100|18193_ ;
  assign \new_Sorter100|18294_  = \new_Sorter100|18194_  & \new_Sorter100|18195_ ;
  assign \new_Sorter100|18295_  = \new_Sorter100|18194_  | \new_Sorter100|18195_ ;
  assign \new_Sorter100|18296_  = \new_Sorter100|18196_  & \new_Sorter100|18197_ ;
  assign \new_Sorter100|18297_  = \new_Sorter100|18196_  | \new_Sorter100|18197_ ;
  assign \new_Sorter100|18298_  = \new_Sorter100|18198_  & \new_Sorter100|18199_ ;
  assign \new_Sorter100|18299_  = \new_Sorter100|18198_  | \new_Sorter100|18199_ ;
  assign \new_Sorter100|18300_  = \new_Sorter100|18200_ ;
  assign \new_Sorter100|18399_  = \new_Sorter100|18299_ ;
  assign \new_Sorter100|18301_  = \new_Sorter100|18201_  & \new_Sorter100|18202_ ;
  assign \new_Sorter100|18302_  = \new_Sorter100|18201_  | \new_Sorter100|18202_ ;
  assign \new_Sorter100|18303_  = \new_Sorter100|18203_  & \new_Sorter100|18204_ ;
  assign \new_Sorter100|18304_  = \new_Sorter100|18203_  | \new_Sorter100|18204_ ;
  assign \new_Sorter100|18305_  = \new_Sorter100|18205_  & \new_Sorter100|18206_ ;
  assign \new_Sorter100|18306_  = \new_Sorter100|18205_  | \new_Sorter100|18206_ ;
  assign \new_Sorter100|18307_  = \new_Sorter100|18207_  & \new_Sorter100|18208_ ;
  assign \new_Sorter100|18308_  = \new_Sorter100|18207_  | \new_Sorter100|18208_ ;
  assign \new_Sorter100|18309_  = \new_Sorter100|18209_  & \new_Sorter100|18210_ ;
  assign \new_Sorter100|18310_  = \new_Sorter100|18209_  | \new_Sorter100|18210_ ;
  assign \new_Sorter100|18311_  = \new_Sorter100|18211_  & \new_Sorter100|18212_ ;
  assign \new_Sorter100|18312_  = \new_Sorter100|18211_  | \new_Sorter100|18212_ ;
  assign \new_Sorter100|18313_  = \new_Sorter100|18213_  & \new_Sorter100|18214_ ;
  assign \new_Sorter100|18314_  = \new_Sorter100|18213_  | \new_Sorter100|18214_ ;
  assign \new_Sorter100|18315_  = \new_Sorter100|18215_  & \new_Sorter100|18216_ ;
  assign \new_Sorter100|18316_  = \new_Sorter100|18215_  | \new_Sorter100|18216_ ;
  assign \new_Sorter100|18317_  = \new_Sorter100|18217_  & \new_Sorter100|18218_ ;
  assign \new_Sorter100|18318_  = \new_Sorter100|18217_  | \new_Sorter100|18218_ ;
  assign \new_Sorter100|18319_  = \new_Sorter100|18219_  & \new_Sorter100|18220_ ;
  assign \new_Sorter100|18320_  = \new_Sorter100|18219_  | \new_Sorter100|18220_ ;
  assign \new_Sorter100|18321_  = \new_Sorter100|18221_  & \new_Sorter100|18222_ ;
  assign \new_Sorter100|18322_  = \new_Sorter100|18221_  | \new_Sorter100|18222_ ;
  assign \new_Sorter100|18323_  = \new_Sorter100|18223_  & \new_Sorter100|18224_ ;
  assign \new_Sorter100|18324_  = \new_Sorter100|18223_  | \new_Sorter100|18224_ ;
  assign \new_Sorter100|18325_  = \new_Sorter100|18225_  & \new_Sorter100|18226_ ;
  assign \new_Sorter100|18326_  = \new_Sorter100|18225_  | \new_Sorter100|18226_ ;
  assign \new_Sorter100|18327_  = \new_Sorter100|18227_  & \new_Sorter100|18228_ ;
  assign \new_Sorter100|18328_  = \new_Sorter100|18227_  | \new_Sorter100|18228_ ;
  assign \new_Sorter100|18329_  = \new_Sorter100|18229_  & \new_Sorter100|18230_ ;
  assign \new_Sorter100|18330_  = \new_Sorter100|18229_  | \new_Sorter100|18230_ ;
  assign \new_Sorter100|18331_  = \new_Sorter100|18231_  & \new_Sorter100|18232_ ;
  assign \new_Sorter100|18332_  = \new_Sorter100|18231_  | \new_Sorter100|18232_ ;
  assign \new_Sorter100|18333_  = \new_Sorter100|18233_  & \new_Sorter100|18234_ ;
  assign \new_Sorter100|18334_  = \new_Sorter100|18233_  | \new_Sorter100|18234_ ;
  assign \new_Sorter100|18335_  = \new_Sorter100|18235_  & \new_Sorter100|18236_ ;
  assign \new_Sorter100|18336_  = \new_Sorter100|18235_  | \new_Sorter100|18236_ ;
  assign \new_Sorter100|18337_  = \new_Sorter100|18237_  & \new_Sorter100|18238_ ;
  assign \new_Sorter100|18338_  = \new_Sorter100|18237_  | \new_Sorter100|18238_ ;
  assign \new_Sorter100|18339_  = \new_Sorter100|18239_  & \new_Sorter100|18240_ ;
  assign \new_Sorter100|18340_  = \new_Sorter100|18239_  | \new_Sorter100|18240_ ;
  assign \new_Sorter100|18341_  = \new_Sorter100|18241_  & \new_Sorter100|18242_ ;
  assign \new_Sorter100|18342_  = \new_Sorter100|18241_  | \new_Sorter100|18242_ ;
  assign \new_Sorter100|18343_  = \new_Sorter100|18243_  & \new_Sorter100|18244_ ;
  assign \new_Sorter100|18344_  = \new_Sorter100|18243_  | \new_Sorter100|18244_ ;
  assign \new_Sorter100|18345_  = \new_Sorter100|18245_  & \new_Sorter100|18246_ ;
  assign \new_Sorter100|18346_  = \new_Sorter100|18245_  | \new_Sorter100|18246_ ;
  assign \new_Sorter100|18347_  = \new_Sorter100|18247_  & \new_Sorter100|18248_ ;
  assign \new_Sorter100|18348_  = \new_Sorter100|18247_  | \new_Sorter100|18248_ ;
  assign \new_Sorter100|18349_  = \new_Sorter100|18249_  & \new_Sorter100|18250_ ;
  assign \new_Sorter100|18350_  = \new_Sorter100|18249_  | \new_Sorter100|18250_ ;
  assign \new_Sorter100|18351_  = \new_Sorter100|18251_  & \new_Sorter100|18252_ ;
  assign \new_Sorter100|18352_  = \new_Sorter100|18251_  | \new_Sorter100|18252_ ;
  assign \new_Sorter100|18353_  = \new_Sorter100|18253_  & \new_Sorter100|18254_ ;
  assign \new_Sorter100|18354_  = \new_Sorter100|18253_  | \new_Sorter100|18254_ ;
  assign \new_Sorter100|18355_  = \new_Sorter100|18255_  & \new_Sorter100|18256_ ;
  assign \new_Sorter100|18356_  = \new_Sorter100|18255_  | \new_Sorter100|18256_ ;
  assign \new_Sorter100|18357_  = \new_Sorter100|18257_  & \new_Sorter100|18258_ ;
  assign \new_Sorter100|18358_  = \new_Sorter100|18257_  | \new_Sorter100|18258_ ;
  assign \new_Sorter100|18359_  = \new_Sorter100|18259_  & \new_Sorter100|18260_ ;
  assign \new_Sorter100|18360_  = \new_Sorter100|18259_  | \new_Sorter100|18260_ ;
  assign \new_Sorter100|18361_  = \new_Sorter100|18261_  & \new_Sorter100|18262_ ;
  assign \new_Sorter100|18362_  = \new_Sorter100|18261_  | \new_Sorter100|18262_ ;
  assign \new_Sorter100|18363_  = \new_Sorter100|18263_  & \new_Sorter100|18264_ ;
  assign \new_Sorter100|18364_  = \new_Sorter100|18263_  | \new_Sorter100|18264_ ;
  assign \new_Sorter100|18365_  = \new_Sorter100|18265_  & \new_Sorter100|18266_ ;
  assign \new_Sorter100|18366_  = \new_Sorter100|18265_  | \new_Sorter100|18266_ ;
  assign \new_Sorter100|18367_  = \new_Sorter100|18267_  & \new_Sorter100|18268_ ;
  assign \new_Sorter100|18368_  = \new_Sorter100|18267_  | \new_Sorter100|18268_ ;
  assign \new_Sorter100|18369_  = \new_Sorter100|18269_  & \new_Sorter100|18270_ ;
  assign \new_Sorter100|18370_  = \new_Sorter100|18269_  | \new_Sorter100|18270_ ;
  assign \new_Sorter100|18371_  = \new_Sorter100|18271_  & \new_Sorter100|18272_ ;
  assign \new_Sorter100|18372_  = \new_Sorter100|18271_  | \new_Sorter100|18272_ ;
  assign \new_Sorter100|18373_  = \new_Sorter100|18273_  & \new_Sorter100|18274_ ;
  assign \new_Sorter100|18374_  = \new_Sorter100|18273_  | \new_Sorter100|18274_ ;
  assign \new_Sorter100|18375_  = \new_Sorter100|18275_  & \new_Sorter100|18276_ ;
  assign \new_Sorter100|18376_  = \new_Sorter100|18275_  | \new_Sorter100|18276_ ;
  assign \new_Sorter100|18377_  = \new_Sorter100|18277_  & \new_Sorter100|18278_ ;
  assign \new_Sorter100|18378_  = \new_Sorter100|18277_  | \new_Sorter100|18278_ ;
  assign \new_Sorter100|18379_  = \new_Sorter100|18279_  & \new_Sorter100|18280_ ;
  assign \new_Sorter100|18380_  = \new_Sorter100|18279_  | \new_Sorter100|18280_ ;
  assign \new_Sorter100|18381_  = \new_Sorter100|18281_  & \new_Sorter100|18282_ ;
  assign \new_Sorter100|18382_  = \new_Sorter100|18281_  | \new_Sorter100|18282_ ;
  assign \new_Sorter100|18383_  = \new_Sorter100|18283_  & \new_Sorter100|18284_ ;
  assign \new_Sorter100|18384_  = \new_Sorter100|18283_  | \new_Sorter100|18284_ ;
  assign \new_Sorter100|18385_  = \new_Sorter100|18285_  & \new_Sorter100|18286_ ;
  assign \new_Sorter100|18386_  = \new_Sorter100|18285_  | \new_Sorter100|18286_ ;
  assign \new_Sorter100|18387_  = \new_Sorter100|18287_  & \new_Sorter100|18288_ ;
  assign \new_Sorter100|18388_  = \new_Sorter100|18287_  | \new_Sorter100|18288_ ;
  assign \new_Sorter100|18389_  = \new_Sorter100|18289_  & \new_Sorter100|18290_ ;
  assign \new_Sorter100|18390_  = \new_Sorter100|18289_  | \new_Sorter100|18290_ ;
  assign \new_Sorter100|18391_  = \new_Sorter100|18291_  & \new_Sorter100|18292_ ;
  assign \new_Sorter100|18392_  = \new_Sorter100|18291_  | \new_Sorter100|18292_ ;
  assign \new_Sorter100|18393_  = \new_Sorter100|18293_  & \new_Sorter100|18294_ ;
  assign \new_Sorter100|18394_  = \new_Sorter100|18293_  | \new_Sorter100|18294_ ;
  assign \new_Sorter100|18395_  = \new_Sorter100|18295_  & \new_Sorter100|18296_ ;
  assign \new_Sorter100|18396_  = \new_Sorter100|18295_  | \new_Sorter100|18296_ ;
  assign \new_Sorter100|18397_  = \new_Sorter100|18297_  & \new_Sorter100|18298_ ;
  assign \new_Sorter100|18398_  = \new_Sorter100|18297_  | \new_Sorter100|18298_ ;
  assign \new_Sorter100|18400_  = \new_Sorter100|18300_  & \new_Sorter100|18301_ ;
  assign \new_Sorter100|18401_  = \new_Sorter100|18300_  | \new_Sorter100|18301_ ;
  assign \new_Sorter100|18402_  = \new_Sorter100|18302_  & \new_Sorter100|18303_ ;
  assign \new_Sorter100|18403_  = \new_Sorter100|18302_  | \new_Sorter100|18303_ ;
  assign \new_Sorter100|18404_  = \new_Sorter100|18304_  & \new_Sorter100|18305_ ;
  assign \new_Sorter100|18405_  = \new_Sorter100|18304_  | \new_Sorter100|18305_ ;
  assign \new_Sorter100|18406_  = \new_Sorter100|18306_  & \new_Sorter100|18307_ ;
  assign \new_Sorter100|18407_  = \new_Sorter100|18306_  | \new_Sorter100|18307_ ;
  assign \new_Sorter100|18408_  = \new_Sorter100|18308_  & \new_Sorter100|18309_ ;
  assign \new_Sorter100|18409_  = \new_Sorter100|18308_  | \new_Sorter100|18309_ ;
  assign \new_Sorter100|18410_  = \new_Sorter100|18310_  & \new_Sorter100|18311_ ;
  assign \new_Sorter100|18411_  = \new_Sorter100|18310_  | \new_Sorter100|18311_ ;
  assign \new_Sorter100|18412_  = \new_Sorter100|18312_  & \new_Sorter100|18313_ ;
  assign \new_Sorter100|18413_  = \new_Sorter100|18312_  | \new_Sorter100|18313_ ;
  assign \new_Sorter100|18414_  = \new_Sorter100|18314_  & \new_Sorter100|18315_ ;
  assign \new_Sorter100|18415_  = \new_Sorter100|18314_  | \new_Sorter100|18315_ ;
  assign \new_Sorter100|18416_  = \new_Sorter100|18316_  & \new_Sorter100|18317_ ;
  assign \new_Sorter100|18417_  = \new_Sorter100|18316_  | \new_Sorter100|18317_ ;
  assign \new_Sorter100|18418_  = \new_Sorter100|18318_  & \new_Sorter100|18319_ ;
  assign \new_Sorter100|18419_  = \new_Sorter100|18318_  | \new_Sorter100|18319_ ;
  assign \new_Sorter100|18420_  = \new_Sorter100|18320_  & \new_Sorter100|18321_ ;
  assign \new_Sorter100|18421_  = \new_Sorter100|18320_  | \new_Sorter100|18321_ ;
  assign \new_Sorter100|18422_  = \new_Sorter100|18322_  & \new_Sorter100|18323_ ;
  assign \new_Sorter100|18423_  = \new_Sorter100|18322_  | \new_Sorter100|18323_ ;
  assign \new_Sorter100|18424_  = \new_Sorter100|18324_  & \new_Sorter100|18325_ ;
  assign \new_Sorter100|18425_  = \new_Sorter100|18324_  | \new_Sorter100|18325_ ;
  assign \new_Sorter100|18426_  = \new_Sorter100|18326_  & \new_Sorter100|18327_ ;
  assign \new_Sorter100|18427_  = \new_Sorter100|18326_  | \new_Sorter100|18327_ ;
  assign \new_Sorter100|18428_  = \new_Sorter100|18328_  & \new_Sorter100|18329_ ;
  assign \new_Sorter100|18429_  = \new_Sorter100|18328_  | \new_Sorter100|18329_ ;
  assign \new_Sorter100|18430_  = \new_Sorter100|18330_  & \new_Sorter100|18331_ ;
  assign \new_Sorter100|18431_  = \new_Sorter100|18330_  | \new_Sorter100|18331_ ;
  assign \new_Sorter100|18432_  = \new_Sorter100|18332_  & \new_Sorter100|18333_ ;
  assign \new_Sorter100|18433_  = \new_Sorter100|18332_  | \new_Sorter100|18333_ ;
  assign \new_Sorter100|18434_  = \new_Sorter100|18334_  & \new_Sorter100|18335_ ;
  assign \new_Sorter100|18435_  = \new_Sorter100|18334_  | \new_Sorter100|18335_ ;
  assign \new_Sorter100|18436_  = \new_Sorter100|18336_  & \new_Sorter100|18337_ ;
  assign \new_Sorter100|18437_  = \new_Sorter100|18336_  | \new_Sorter100|18337_ ;
  assign \new_Sorter100|18438_  = \new_Sorter100|18338_  & \new_Sorter100|18339_ ;
  assign \new_Sorter100|18439_  = \new_Sorter100|18338_  | \new_Sorter100|18339_ ;
  assign \new_Sorter100|18440_  = \new_Sorter100|18340_  & \new_Sorter100|18341_ ;
  assign \new_Sorter100|18441_  = \new_Sorter100|18340_  | \new_Sorter100|18341_ ;
  assign \new_Sorter100|18442_  = \new_Sorter100|18342_  & \new_Sorter100|18343_ ;
  assign \new_Sorter100|18443_  = \new_Sorter100|18342_  | \new_Sorter100|18343_ ;
  assign \new_Sorter100|18444_  = \new_Sorter100|18344_  & \new_Sorter100|18345_ ;
  assign \new_Sorter100|18445_  = \new_Sorter100|18344_  | \new_Sorter100|18345_ ;
  assign \new_Sorter100|18446_  = \new_Sorter100|18346_  & \new_Sorter100|18347_ ;
  assign \new_Sorter100|18447_  = \new_Sorter100|18346_  | \new_Sorter100|18347_ ;
  assign \new_Sorter100|18448_  = \new_Sorter100|18348_  & \new_Sorter100|18349_ ;
  assign \new_Sorter100|18449_  = \new_Sorter100|18348_  | \new_Sorter100|18349_ ;
  assign \new_Sorter100|18450_  = \new_Sorter100|18350_  & \new_Sorter100|18351_ ;
  assign \new_Sorter100|18451_  = \new_Sorter100|18350_  | \new_Sorter100|18351_ ;
  assign \new_Sorter100|18452_  = \new_Sorter100|18352_  & \new_Sorter100|18353_ ;
  assign \new_Sorter100|18453_  = \new_Sorter100|18352_  | \new_Sorter100|18353_ ;
  assign \new_Sorter100|18454_  = \new_Sorter100|18354_  & \new_Sorter100|18355_ ;
  assign \new_Sorter100|18455_  = \new_Sorter100|18354_  | \new_Sorter100|18355_ ;
  assign \new_Sorter100|18456_  = \new_Sorter100|18356_  & \new_Sorter100|18357_ ;
  assign \new_Sorter100|18457_  = \new_Sorter100|18356_  | \new_Sorter100|18357_ ;
  assign \new_Sorter100|18458_  = \new_Sorter100|18358_  & \new_Sorter100|18359_ ;
  assign \new_Sorter100|18459_  = \new_Sorter100|18358_  | \new_Sorter100|18359_ ;
  assign \new_Sorter100|18460_  = \new_Sorter100|18360_  & \new_Sorter100|18361_ ;
  assign \new_Sorter100|18461_  = \new_Sorter100|18360_  | \new_Sorter100|18361_ ;
  assign \new_Sorter100|18462_  = \new_Sorter100|18362_  & \new_Sorter100|18363_ ;
  assign \new_Sorter100|18463_  = \new_Sorter100|18362_  | \new_Sorter100|18363_ ;
  assign \new_Sorter100|18464_  = \new_Sorter100|18364_  & \new_Sorter100|18365_ ;
  assign \new_Sorter100|18465_  = \new_Sorter100|18364_  | \new_Sorter100|18365_ ;
  assign \new_Sorter100|18466_  = \new_Sorter100|18366_  & \new_Sorter100|18367_ ;
  assign \new_Sorter100|18467_  = \new_Sorter100|18366_  | \new_Sorter100|18367_ ;
  assign \new_Sorter100|18468_  = \new_Sorter100|18368_  & \new_Sorter100|18369_ ;
  assign \new_Sorter100|18469_  = \new_Sorter100|18368_  | \new_Sorter100|18369_ ;
  assign \new_Sorter100|18470_  = \new_Sorter100|18370_  & \new_Sorter100|18371_ ;
  assign \new_Sorter100|18471_  = \new_Sorter100|18370_  | \new_Sorter100|18371_ ;
  assign \new_Sorter100|18472_  = \new_Sorter100|18372_  & \new_Sorter100|18373_ ;
  assign \new_Sorter100|18473_  = \new_Sorter100|18372_  | \new_Sorter100|18373_ ;
  assign \new_Sorter100|18474_  = \new_Sorter100|18374_  & \new_Sorter100|18375_ ;
  assign \new_Sorter100|18475_  = \new_Sorter100|18374_  | \new_Sorter100|18375_ ;
  assign \new_Sorter100|18476_  = \new_Sorter100|18376_  & \new_Sorter100|18377_ ;
  assign \new_Sorter100|18477_  = \new_Sorter100|18376_  | \new_Sorter100|18377_ ;
  assign \new_Sorter100|18478_  = \new_Sorter100|18378_  & \new_Sorter100|18379_ ;
  assign \new_Sorter100|18479_  = \new_Sorter100|18378_  | \new_Sorter100|18379_ ;
  assign \new_Sorter100|18480_  = \new_Sorter100|18380_  & \new_Sorter100|18381_ ;
  assign \new_Sorter100|18481_  = \new_Sorter100|18380_  | \new_Sorter100|18381_ ;
  assign \new_Sorter100|18482_  = \new_Sorter100|18382_  & \new_Sorter100|18383_ ;
  assign \new_Sorter100|18483_  = \new_Sorter100|18382_  | \new_Sorter100|18383_ ;
  assign \new_Sorter100|18484_  = \new_Sorter100|18384_  & \new_Sorter100|18385_ ;
  assign \new_Sorter100|18485_  = \new_Sorter100|18384_  | \new_Sorter100|18385_ ;
  assign \new_Sorter100|18486_  = \new_Sorter100|18386_  & \new_Sorter100|18387_ ;
  assign \new_Sorter100|18487_  = \new_Sorter100|18386_  | \new_Sorter100|18387_ ;
  assign \new_Sorter100|18488_  = \new_Sorter100|18388_  & \new_Sorter100|18389_ ;
  assign \new_Sorter100|18489_  = \new_Sorter100|18388_  | \new_Sorter100|18389_ ;
  assign \new_Sorter100|18490_  = \new_Sorter100|18390_  & \new_Sorter100|18391_ ;
  assign \new_Sorter100|18491_  = \new_Sorter100|18390_  | \new_Sorter100|18391_ ;
  assign \new_Sorter100|18492_  = \new_Sorter100|18392_  & \new_Sorter100|18393_ ;
  assign \new_Sorter100|18493_  = \new_Sorter100|18392_  | \new_Sorter100|18393_ ;
  assign \new_Sorter100|18494_  = \new_Sorter100|18394_  & \new_Sorter100|18395_ ;
  assign \new_Sorter100|18495_  = \new_Sorter100|18394_  | \new_Sorter100|18395_ ;
  assign \new_Sorter100|18496_  = \new_Sorter100|18396_  & \new_Sorter100|18397_ ;
  assign \new_Sorter100|18497_  = \new_Sorter100|18396_  | \new_Sorter100|18397_ ;
  assign \new_Sorter100|18498_  = \new_Sorter100|18398_  & \new_Sorter100|18399_ ;
  assign \new_Sorter100|18499_  = \new_Sorter100|18398_  | \new_Sorter100|18399_ ;
  assign \new_Sorter100|18500_  = \new_Sorter100|18400_ ;
  assign \new_Sorter100|18599_  = \new_Sorter100|18499_ ;
  assign \new_Sorter100|18501_  = \new_Sorter100|18401_  & \new_Sorter100|18402_ ;
  assign \new_Sorter100|18502_  = \new_Sorter100|18401_  | \new_Sorter100|18402_ ;
  assign \new_Sorter100|18503_  = \new_Sorter100|18403_  & \new_Sorter100|18404_ ;
  assign \new_Sorter100|18504_  = \new_Sorter100|18403_  | \new_Sorter100|18404_ ;
  assign \new_Sorter100|18505_  = \new_Sorter100|18405_  & \new_Sorter100|18406_ ;
  assign \new_Sorter100|18506_  = \new_Sorter100|18405_  | \new_Sorter100|18406_ ;
  assign \new_Sorter100|18507_  = \new_Sorter100|18407_  & \new_Sorter100|18408_ ;
  assign \new_Sorter100|18508_  = \new_Sorter100|18407_  | \new_Sorter100|18408_ ;
  assign \new_Sorter100|18509_  = \new_Sorter100|18409_  & \new_Sorter100|18410_ ;
  assign \new_Sorter100|18510_  = \new_Sorter100|18409_  | \new_Sorter100|18410_ ;
  assign \new_Sorter100|18511_  = \new_Sorter100|18411_  & \new_Sorter100|18412_ ;
  assign \new_Sorter100|18512_  = \new_Sorter100|18411_  | \new_Sorter100|18412_ ;
  assign \new_Sorter100|18513_  = \new_Sorter100|18413_  & \new_Sorter100|18414_ ;
  assign \new_Sorter100|18514_  = \new_Sorter100|18413_  | \new_Sorter100|18414_ ;
  assign \new_Sorter100|18515_  = \new_Sorter100|18415_  & \new_Sorter100|18416_ ;
  assign \new_Sorter100|18516_  = \new_Sorter100|18415_  | \new_Sorter100|18416_ ;
  assign \new_Sorter100|18517_  = \new_Sorter100|18417_  & \new_Sorter100|18418_ ;
  assign \new_Sorter100|18518_  = \new_Sorter100|18417_  | \new_Sorter100|18418_ ;
  assign \new_Sorter100|18519_  = \new_Sorter100|18419_  & \new_Sorter100|18420_ ;
  assign \new_Sorter100|18520_  = \new_Sorter100|18419_  | \new_Sorter100|18420_ ;
  assign \new_Sorter100|18521_  = \new_Sorter100|18421_  & \new_Sorter100|18422_ ;
  assign \new_Sorter100|18522_  = \new_Sorter100|18421_  | \new_Sorter100|18422_ ;
  assign \new_Sorter100|18523_  = \new_Sorter100|18423_  & \new_Sorter100|18424_ ;
  assign \new_Sorter100|18524_  = \new_Sorter100|18423_  | \new_Sorter100|18424_ ;
  assign \new_Sorter100|18525_  = \new_Sorter100|18425_  & \new_Sorter100|18426_ ;
  assign \new_Sorter100|18526_  = \new_Sorter100|18425_  | \new_Sorter100|18426_ ;
  assign \new_Sorter100|18527_  = \new_Sorter100|18427_  & \new_Sorter100|18428_ ;
  assign \new_Sorter100|18528_  = \new_Sorter100|18427_  | \new_Sorter100|18428_ ;
  assign \new_Sorter100|18529_  = \new_Sorter100|18429_  & \new_Sorter100|18430_ ;
  assign \new_Sorter100|18530_  = \new_Sorter100|18429_  | \new_Sorter100|18430_ ;
  assign \new_Sorter100|18531_  = \new_Sorter100|18431_  & \new_Sorter100|18432_ ;
  assign \new_Sorter100|18532_  = \new_Sorter100|18431_  | \new_Sorter100|18432_ ;
  assign \new_Sorter100|18533_  = \new_Sorter100|18433_  & \new_Sorter100|18434_ ;
  assign \new_Sorter100|18534_  = \new_Sorter100|18433_  | \new_Sorter100|18434_ ;
  assign \new_Sorter100|18535_  = \new_Sorter100|18435_  & \new_Sorter100|18436_ ;
  assign \new_Sorter100|18536_  = \new_Sorter100|18435_  | \new_Sorter100|18436_ ;
  assign \new_Sorter100|18537_  = \new_Sorter100|18437_  & \new_Sorter100|18438_ ;
  assign \new_Sorter100|18538_  = \new_Sorter100|18437_  | \new_Sorter100|18438_ ;
  assign \new_Sorter100|18539_  = \new_Sorter100|18439_  & \new_Sorter100|18440_ ;
  assign \new_Sorter100|18540_  = \new_Sorter100|18439_  | \new_Sorter100|18440_ ;
  assign \new_Sorter100|18541_  = \new_Sorter100|18441_  & \new_Sorter100|18442_ ;
  assign \new_Sorter100|18542_  = \new_Sorter100|18441_  | \new_Sorter100|18442_ ;
  assign \new_Sorter100|18543_  = \new_Sorter100|18443_  & \new_Sorter100|18444_ ;
  assign \new_Sorter100|18544_  = \new_Sorter100|18443_  | \new_Sorter100|18444_ ;
  assign \new_Sorter100|18545_  = \new_Sorter100|18445_  & \new_Sorter100|18446_ ;
  assign \new_Sorter100|18546_  = \new_Sorter100|18445_  | \new_Sorter100|18446_ ;
  assign \new_Sorter100|18547_  = \new_Sorter100|18447_  & \new_Sorter100|18448_ ;
  assign \new_Sorter100|18548_  = \new_Sorter100|18447_  | \new_Sorter100|18448_ ;
  assign \new_Sorter100|18549_  = \new_Sorter100|18449_  & \new_Sorter100|18450_ ;
  assign \new_Sorter100|18550_  = \new_Sorter100|18449_  | \new_Sorter100|18450_ ;
  assign \new_Sorter100|18551_  = \new_Sorter100|18451_  & \new_Sorter100|18452_ ;
  assign \new_Sorter100|18552_  = \new_Sorter100|18451_  | \new_Sorter100|18452_ ;
  assign \new_Sorter100|18553_  = \new_Sorter100|18453_  & \new_Sorter100|18454_ ;
  assign \new_Sorter100|18554_  = \new_Sorter100|18453_  | \new_Sorter100|18454_ ;
  assign \new_Sorter100|18555_  = \new_Sorter100|18455_  & \new_Sorter100|18456_ ;
  assign \new_Sorter100|18556_  = \new_Sorter100|18455_  | \new_Sorter100|18456_ ;
  assign \new_Sorter100|18557_  = \new_Sorter100|18457_  & \new_Sorter100|18458_ ;
  assign \new_Sorter100|18558_  = \new_Sorter100|18457_  | \new_Sorter100|18458_ ;
  assign \new_Sorter100|18559_  = \new_Sorter100|18459_  & \new_Sorter100|18460_ ;
  assign \new_Sorter100|18560_  = \new_Sorter100|18459_  | \new_Sorter100|18460_ ;
  assign \new_Sorter100|18561_  = \new_Sorter100|18461_  & \new_Sorter100|18462_ ;
  assign \new_Sorter100|18562_  = \new_Sorter100|18461_  | \new_Sorter100|18462_ ;
  assign \new_Sorter100|18563_  = \new_Sorter100|18463_  & \new_Sorter100|18464_ ;
  assign \new_Sorter100|18564_  = \new_Sorter100|18463_  | \new_Sorter100|18464_ ;
  assign \new_Sorter100|18565_  = \new_Sorter100|18465_  & \new_Sorter100|18466_ ;
  assign \new_Sorter100|18566_  = \new_Sorter100|18465_  | \new_Sorter100|18466_ ;
  assign \new_Sorter100|18567_  = \new_Sorter100|18467_  & \new_Sorter100|18468_ ;
  assign \new_Sorter100|18568_  = \new_Sorter100|18467_  | \new_Sorter100|18468_ ;
  assign \new_Sorter100|18569_  = \new_Sorter100|18469_  & \new_Sorter100|18470_ ;
  assign \new_Sorter100|18570_  = \new_Sorter100|18469_  | \new_Sorter100|18470_ ;
  assign \new_Sorter100|18571_  = \new_Sorter100|18471_  & \new_Sorter100|18472_ ;
  assign \new_Sorter100|18572_  = \new_Sorter100|18471_  | \new_Sorter100|18472_ ;
  assign \new_Sorter100|18573_  = \new_Sorter100|18473_  & \new_Sorter100|18474_ ;
  assign \new_Sorter100|18574_  = \new_Sorter100|18473_  | \new_Sorter100|18474_ ;
  assign \new_Sorter100|18575_  = \new_Sorter100|18475_  & \new_Sorter100|18476_ ;
  assign \new_Sorter100|18576_  = \new_Sorter100|18475_  | \new_Sorter100|18476_ ;
  assign \new_Sorter100|18577_  = \new_Sorter100|18477_  & \new_Sorter100|18478_ ;
  assign \new_Sorter100|18578_  = \new_Sorter100|18477_  | \new_Sorter100|18478_ ;
  assign \new_Sorter100|18579_  = \new_Sorter100|18479_  & \new_Sorter100|18480_ ;
  assign \new_Sorter100|18580_  = \new_Sorter100|18479_  | \new_Sorter100|18480_ ;
  assign \new_Sorter100|18581_  = \new_Sorter100|18481_  & \new_Sorter100|18482_ ;
  assign \new_Sorter100|18582_  = \new_Sorter100|18481_  | \new_Sorter100|18482_ ;
  assign \new_Sorter100|18583_  = \new_Sorter100|18483_  & \new_Sorter100|18484_ ;
  assign \new_Sorter100|18584_  = \new_Sorter100|18483_  | \new_Sorter100|18484_ ;
  assign \new_Sorter100|18585_  = \new_Sorter100|18485_  & \new_Sorter100|18486_ ;
  assign \new_Sorter100|18586_  = \new_Sorter100|18485_  | \new_Sorter100|18486_ ;
  assign \new_Sorter100|18587_  = \new_Sorter100|18487_  & \new_Sorter100|18488_ ;
  assign \new_Sorter100|18588_  = \new_Sorter100|18487_  | \new_Sorter100|18488_ ;
  assign \new_Sorter100|18589_  = \new_Sorter100|18489_  & \new_Sorter100|18490_ ;
  assign \new_Sorter100|18590_  = \new_Sorter100|18489_  | \new_Sorter100|18490_ ;
  assign \new_Sorter100|18591_  = \new_Sorter100|18491_  & \new_Sorter100|18492_ ;
  assign \new_Sorter100|18592_  = \new_Sorter100|18491_  | \new_Sorter100|18492_ ;
  assign \new_Sorter100|18593_  = \new_Sorter100|18493_  & \new_Sorter100|18494_ ;
  assign \new_Sorter100|18594_  = \new_Sorter100|18493_  | \new_Sorter100|18494_ ;
  assign \new_Sorter100|18595_  = \new_Sorter100|18495_  & \new_Sorter100|18496_ ;
  assign \new_Sorter100|18596_  = \new_Sorter100|18495_  | \new_Sorter100|18496_ ;
  assign \new_Sorter100|18597_  = \new_Sorter100|18497_  & \new_Sorter100|18498_ ;
  assign \new_Sorter100|18598_  = \new_Sorter100|18497_  | \new_Sorter100|18498_ ;
  assign \new_Sorter100|18600_  = \new_Sorter100|18500_  & \new_Sorter100|18501_ ;
  assign \new_Sorter100|18601_  = \new_Sorter100|18500_  | \new_Sorter100|18501_ ;
  assign \new_Sorter100|18602_  = \new_Sorter100|18502_  & \new_Sorter100|18503_ ;
  assign \new_Sorter100|18603_  = \new_Sorter100|18502_  | \new_Sorter100|18503_ ;
  assign \new_Sorter100|18604_  = \new_Sorter100|18504_  & \new_Sorter100|18505_ ;
  assign \new_Sorter100|18605_  = \new_Sorter100|18504_  | \new_Sorter100|18505_ ;
  assign \new_Sorter100|18606_  = \new_Sorter100|18506_  & \new_Sorter100|18507_ ;
  assign \new_Sorter100|18607_  = \new_Sorter100|18506_  | \new_Sorter100|18507_ ;
  assign \new_Sorter100|18608_  = \new_Sorter100|18508_  & \new_Sorter100|18509_ ;
  assign \new_Sorter100|18609_  = \new_Sorter100|18508_  | \new_Sorter100|18509_ ;
  assign \new_Sorter100|18610_  = \new_Sorter100|18510_  & \new_Sorter100|18511_ ;
  assign \new_Sorter100|18611_  = \new_Sorter100|18510_  | \new_Sorter100|18511_ ;
  assign \new_Sorter100|18612_  = \new_Sorter100|18512_  & \new_Sorter100|18513_ ;
  assign \new_Sorter100|18613_  = \new_Sorter100|18512_  | \new_Sorter100|18513_ ;
  assign \new_Sorter100|18614_  = \new_Sorter100|18514_  & \new_Sorter100|18515_ ;
  assign \new_Sorter100|18615_  = \new_Sorter100|18514_  | \new_Sorter100|18515_ ;
  assign \new_Sorter100|18616_  = \new_Sorter100|18516_  & \new_Sorter100|18517_ ;
  assign \new_Sorter100|18617_  = \new_Sorter100|18516_  | \new_Sorter100|18517_ ;
  assign \new_Sorter100|18618_  = \new_Sorter100|18518_  & \new_Sorter100|18519_ ;
  assign \new_Sorter100|18619_  = \new_Sorter100|18518_  | \new_Sorter100|18519_ ;
  assign \new_Sorter100|18620_  = \new_Sorter100|18520_  & \new_Sorter100|18521_ ;
  assign \new_Sorter100|18621_  = \new_Sorter100|18520_  | \new_Sorter100|18521_ ;
  assign \new_Sorter100|18622_  = \new_Sorter100|18522_  & \new_Sorter100|18523_ ;
  assign \new_Sorter100|18623_  = \new_Sorter100|18522_  | \new_Sorter100|18523_ ;
  assign \new_Sorter100|18624_  = \new_Sorter100|18524_  & \new_Sorter100|18525_ ;
  assign \new_Sorter100|18625_  = \new_Sorter100|18524_  | \new_Sorter100|18525_ ;
  assign \new_Sorter100|18626_  = \new_Sorter100|18526_  & \new_Sorter100|18527_ ;
  assign \new_Sorter100|18627_  = \new_Sorter100|18526_  | \new_Sorter100|18527_ ;
  assign \new_Sorter100|18628_  = \new_Sorter100|18528_  & \new_Sorter100|18529_ ;
  assign \new_Sorter100|18629_  = \new_Sorter100|18528_  | \new_Sorter100|18529_ ;
  assign \new_Sorter100|18630_  = \new_Sorter100|18530_  & \new_Sorter100|18531_ ;
  assign \new_Sorter100|18631_  = \new_Sorter100|18530_  | \new_Sorter100|18531_ ;
  assign \new_Sorter100|18632_  = \new_Sorter100|18532_  & \new_Sorter100|18533_ ;
  assign \new_Sorter100|18633_  = \new_Sorter100|18532_  | \new_Sorter100|18533_ ;
  assign \new_Sorter100|18634_  = \new_Sorter100|18534_  & \new_Sorter100|18535_ ;
  assign \new_Sorter100|18635_  = \new_Sorter100|18534_  | \new_Sorter100|18535_ ;
  assign \new_Sorter100|18636_  = \new_Sorter100|18536_  & \new_Sorter100|18537_ ;
  assign \new_Sorter100|18637_  = \new_Sorter100|18536_  | \new_Sorter100|18537_ ;
  assign \new_Sorter100|18638_  = \new_Sorter100|18538_  & \new_Sorter100|18539_ ;
  assign \new_Sorter100|18639_  = \new_Sorter100|18538_  | \new_Sorter100|18539_ ;
  assign \new_Sorter100|18640_  = \new_Sorter100|18540_  & \new_Sorter100|18541_ ;
  assign \new_Sorter100|18641_  = \new_Sorter100|18540_  | \new_Sorter100|18541_ ;
  assign \new_Sorter100|18642_  = \new_Sorter100|18542_  & \new_Sorter100|18543_ ;
  assign \new_Sorter100|18643_  = \new_Sorter100|18542_  | \new_Sorter100|18543_ ;
  assign \new_Sorter100|18644_  = \new_Sorter100|18544_  & \new_Sorter100|18545_ ;
  assign \new_Sorter100|18645_  = \new_Sorter100|18544_  | \new_Sorter100|18545_ ;
  assign \new_Sorter100|18646_  = \new_Sorter100|18546_  & \new_Sorter100|18547_ ;
  assign \new_Sorter100|18647_  = \new_Sorter100|18546_  | \new_Sorter100|18547_ ;
  assign \new_Sorter100|18648_  = \new_Sorter100|18548_  & \new_Sorter100|18549_ ;
  assign \new_Sorter100|18649_  = \new_Sorter100|18548_  | \new_Sorter100|18549_ ;
  assign \new_Sorter100|18650_  = \new_Sorter100|18550_  & \new_Sorter100|18551_ ;
  assign \new_Sorter100|18651_  = \new_Sorter100|18550_  | \new_Sorter100|18551_ ;
  assign \new_Sorter100|18652_  = \new_Sorter100|18552_  & \new_Sorter100|18553_ ;
  assign \new_Sorter100|18653_  = \new_Sorter100|18552_  | \new_Sorter100|18553_ ;
  assign \new_Sorter100|18654_  = \new_Sorter100|18554_  & \new_Sorter100|18555_ ;
  assign \new_Sorter100|18655_  = \new_Sorter100|18554_  | \new_Sorter100|18555_ ;
  assign \new_Sorter100|18656_  = \new_Sorter100|18556_  & \new_Sorter100|18557_ ;
  assign \new_Sorter100|18657_  = \new_Sorter100|18556_  | \new_Sorter100|18557_ ;
  assign \new_Sorter100|18658_  = \new_Sorter100|18558_  & \new_Sorter100|18559_ ;
  assign \new_Sorter100|18659_  = \new_Sorter100|18558_  | \new_Sorter100|18559_ ;
  assign \new_Sorter100|18660_  = \new_Sorter100|18560_  & \new_Sorter100|18561_ ;
  assign \new_Sorter100|18661_  = \new_Sorter100|18560_  | \new_Sorter100|18561_ ;
  assign \new_Sorter100|18662_  = \new_Sorter100|18562_  & \new_Sorter100|18563_ ;
  assign \new_Sorter100|18663_  = \new_Sorter100|18562_  | \new_Sorter100|18563_ ;
  assign \new_Sorter100|18664_  = \new_Sorter100|18564_  & \new_Sorter100|18565_ ;
  assign \new_Sorter100|18665_  = \new_Sorter100|18564_  | \new_Sorter100|18565_ ;
  assign \new_Sorter100|18666_  = \new_Sorter100|18566_  & \new_Sorter100|18567_ ;
  assign \new_Sorter100|18667_  = \new_Sorter100|18566_  | \new_Sorter100|18567_ ;
  assign \new_Sorter100|18668_  = \new_Sorter100|18568_  & \new_Sorter100|18569_ ;
  assign \new_Sorter100|18669_  = \new_Sorter100|18568_  | \new_Sorter100|18569_ ;
  assign \new_Sorter100|18670_  = \new_Sorter100|18570_  & \new_Sorter100|18571_ ;
  assign \new_Sorter100|18671_  = \new_Sorter100|18570_  | \new_Sorter100|18571_ ;
  assign \new_Sorter100|18672_  = \new_Sorter100|18572_  & \new_Sorter100|18573_ ;
  assign \new_Sorter100|18673_  = \new_Sorter100|18572_  | \new_Sorter100|18573_ ;
  assign \new_Sorter100|18674_  = \new_Sorter100|18574_  & \new_Sorter100|18575_ ;
  assign \new_Sorter100|18675_  = \new_Sorter100|18574_  | \new_Sorter100|18575_ ;
  assign \new_Sorter100|18676_  = \new_Sorter100|18576_  & \new_Sorter100|18577_ ;
  assign \new_Sorter100|18677_  = \new_Sorter100|18576_  | \new_Sorter100|18577_ ;
  assign \new_Sorter100|18678_  = \new_Sorter100|18578_  & \new_Sorter100|18579_ ;
  assign \new_Sorter100|18679_  = \new_Sorter100|18578_  | \new_Sorter100|18579_ ;
  assign \new_Sorter100|18680_  = \new_Sorter100|18580_  & \new_Sorter100|18581_ ;
  assign \new_Sorter100|18681_  = \new_Sorter100|18580_  | \new_Sorter100|18581_ ;
  assign \new_Sorter100|18682_  = \new_Sorter100|18582_  & \new_Sorter100|18583_ ;
  assign \new_Sorter100|18683_  = \new_Sorter100|18582_  | \new_Sorter100|18583_ ;
  assign \new_Sorter100|18684_  = \new_Sorter100|18584_  & \new_Sorter100|18585_ ;
  assign \new_Sorter100|18685_  = \new_Sorter100|18584_  | \new_Sorter100|18585_ ;
  assign \new_Sorter100|18686_  = \new_Sorter100|18586_  & \new_Sorter100|18587_ ;
  assign \new_Sorter100|18687_  = \new_Sorter100|18586_  | \new_Sorter100|18587_ ;
  assign \new_Sorter100|18688_  = \new_Sorter100|18588_  & \new_Sorter100|18589_ ;
  assign \new_Sorter100|18689_  = \new_Sorter100|18588_  | \new_Sorter100|18589_ ;
  assign \new_Sorter100|18690_  = \new_Sorter100|18590_  & \new_Sorter100|18591_ ;
  assign \new_Sorter100|18691_  = \new_Sorter100|18590_  | \new_Sorter100|18591_ ;
  assign \new_Sorter100|18692_  = \new_Sorter100|18592_  & \new_Sorter100|18593_ ;
  assign \new_Sorter100|18693_  = \new_Sorter100|18592_  | \new_Sorter100|18593_ ;
  assign \new_Sorter100|18694_  = \new_Sorter100|18594_  & \new_Sorter100|18595_ ;
  assign \new_Sorter100|18695_  = \new_Sorter100|18594_  | \new_Sorter100|18595_ ;
  assign \new_Sorter100|18696_  = \new_Sorter100|18596_  & \new_Sorter100|18597_ ;
  assign \new_Sorter100|18697_  = \new_Sorter100|18596_  | \new_Sorter100|18597_ ;
  assign \new_Sorter100|18698_  = \new_Sorter100|18598_  & \new_Sorter100|18599_ ;
  assign \new_Sorter100|18699_  = \new_Sorter100|18598_  | \new_Sorter100|18599_ ;
  assign \new_Sorter100|18700_  = \new_Sorter100|18600_ ;
  assign \new_Sorter100|18799_  = \new_Sorter100|18699_ ;
  assign \new_Sorter100|18701_  = \new_Sorter100|18601_  & \new_Sorter100|18602_ ;
  assign \new_Sorter100|18702_  = \new_Sorter100|18601_  | \new_Sorter100|18602_ ;
  assign \new_Sorter100|18703_  = \new_Sorter100|18603_  & \new_Sorter100|18604_ ;
  assign \new_Sorter100|18704_  = \new_Sorter100|18603_  | \new_Sorter100|18604_ ;
  assign \new_Sorter100|18705_  = \new_Sorter100|18605_  & \new_Sorter100|18606_ ;
  assign \new_Sorter100|18706_  = \new_Sorter100|18605_  | \new_Sorter100|18606_ ;
  assign \new_Sorter100|18707_  = \new_Sorter100|18607_  & \new_Sorter100|18608_ ;
  assign \new_Sorter100|18708_  = \new_Sorter100|18607_  | \new_Sorter100|18608_ ;
  assign \new_Sorter100|18709_  = \new_Sorter100|18609_  & \new_Sorter100|18610_ ;
  assign \new_Sorter100|18710_  = \new_Sorter100|18609_  | \new_Sorter100|18610_ ;
  assign \new_Sorter100|18711_  = \new_Sorter100|18611_  & \new_Sorter100|18612_ ;
  assign \new_Sorter100|18712_  = \new_Sorter100|18611_  | \new_Sorter100|18612_ ;
  assign \new_Sorter100|18713_  = \new_Sorter100|18613_  & \new_Sorter100|18614_ ;
  assign \new_Sorter100|18714_  = \new_Sorter100|18613_  | \new_Sorter100|18614_ ;
  assign \new_Sorter100|18715_  = \new_Sorter100|18615_  & \new_Sorter100|18616_ ;
  assign \new_Sorter100|18716_  = \new_Sorter100|18615_  | \new_Sorter100|18616_ ;
  assign \new_Sorter100|18717_  = \new_Sorter100|18617_  & \new_Sorter100|18618_ ;
  assign \new_Sorter100|18718_  = \new_Sorter100|18617_  | \new_Sorter100|18618_ ;
  assign \new_Sorter100|18719_  = \new_Sorter100|18619_  & \new_Sorter100|18620_ ;
  assign \new_Sorter100|18720_  = \new_Sorter100|18619_  | \new_Sorter100|18620_ ;
  assign \new_Sorter100|18721_  = \new_Sorter100|18621_  & \new_Sorter100|18622_ ;
  assign \new_Sorter100|18722_  = \new_Sorter100|18621_  | \new_Sorter100|18622_ ;
  assign \new_Sorter100|18723_  = \new_Sorter100|18623_  & \new_Sorter100|18624_ ;
  assign \new_Sorter100|18724_  = \new_Sorter100|18623_  | \new_Sorter100|18624_ ;
  assign \new_Sorter100|18725_  = \new_Sorter100|18625_  & \new_Sorter100|18626_ ;
  assign \new_Sorter100|18726_  = \new_Sorter100|18625_  | \new_Sorter100|18626_ ;
  assign \new_Sorter100|18727_  = \new_Sorter100|18627_  & \new_Sorter100|18628_ ;
  assign \new_Sorter100|18728_  = \new_Sorter100|18627_  | \new_Sorter100|18628_ ;
  assign \new_Sorter100|18729_  = \new_Sorter100|18629_  & \new_Sorter100|18630_ ;
  assign \new_Sorter100|18730_  = \new_Sorter100|18629_  | \new_Sorter100|18630_ ;
  assign \new_Sorter100|18731_  = \new_Sorter100|18631_  & \new_Sorter100|18632_ ;
  assign \new_Sorter100|18732_  = \new_Sorter100|18631_  | \new_Sorter100|18632_ ;
  assign \new_Sorter100|18733_  = \new_Sorter100|18633_  & \new_Sorter100|18634_ ;
  assign \new_Sorter100|18734_  = \new_Sorter100|18633_  | \new_Sorter100|18634_ ;
  assign \new_Sorter100|18735_  = \new_Sorter100|18635_  & \new_Sorter100|18636_ ;
  assign \new_Sorter100|18736_  = \new_Sorter100|18635_  | \new_Sorter100|18636_ ;
  assign \new_Sorter100|18737_  = \new_Sorter100|18637_  & \new_Sorter100|18638_ ;
  assign \new_Sorter100|18738_  = \new_Sorter100|18637_  | \new_Sorter100|18638_ ;
  assign \new_Sorter100|18739_  = \new_Sorter100|18639_  & \new_Sorter100|18640_ ;
  assign \new_Sorter100|18740_  = \new_Sorter100|18639_  | \new_Sorter100|18640_ ;
  assign \new_Sorter100|18741_  = \new_Sorter100|18641_  & \new_Sorter100|18642_ ;
  assign \new_Sorter100|18742_  = \new_Sorter100|18641_  | \new_Sorter100|18642_ ;
  assign \new_Sorter100|18743_  = \new_Sorter100|18643_  & \new_Sorter100|18644_ ;
  assign \new_Sorter100|18744_  = \new_Sorter100|18643_  | \new_Sorter100|18644_ ;
  assign \new_Sorter100|18745_  = \new_Sorter100|18645_  & \new_Sorter100|18646_ ;
  assign \new_Sorter100|18746_  = \new_Sorter100|18645_  | \new_Sorter100|18646_ ;
  assign \new_Sorter100|18747_  = \new_Sorter100|18647_  & \new_Sorter100|18648_ ;
  assign \new_Sorter100|18748_  = \new_Sorter100|18647_  | \new_Sorter100|18648_ ;
  assign \new_Sorter100|18749_  = \new_Sorter100|18649_  & \new_Sorter100|18650_ ;
  assign \new_Sorter100|18750_  = \new_Sorter100|18649_  | \new_Sorter100|18650_ ;
  assign \new_Sorter100|18751_  = \new_Sorter100|18651_  & \new_Sorter100|18652_ ;
  assign \new_Sorter100|18752_  = \new_Sorter100|18651_  | \new_Sorter100|18652_ ;
  assign \new_Sorter100|18753_  = \new_Sorter100|18653_  & \new_Sorter100|18654_ ;
  assign \new_Sorter100|18754_  = \new_Sorter100|18653_  | \new_Sorter100|18654_ ;
  assign \new_Sorter100|18755_  = \new_Sorter100|18655_  & \new_Sorter100|18656_ ;
  assign \new_Sorter100|18756_  = \new_Sorter100|18655_  | \new_Sorter100|18656_ ;
  assign \new_Sorter100|18757_  = \new_Sorter100|18657_  & \new_Sorter100|18658_ ;
  assign \new_Sorter100|18758_  = \new_Sorter100|18657_  | \new_Sorter100|18658_ ;
  assign \new_Sorter100|18759_  = \new_Sorter100|18659_  & \new_Sorter100|18660_ ;
  assign \new_Sorter100|18760_  = \new_Sorter100|18659_  | \new_Sorter100|18660_ ;
  assign \new_Sorter100|18761_  = \new_Sorter100|18661_  & \new_Sorter100|18662_ ;
  assign \new_Sorter100|18762_  = \new_Sorter100|18661_  | \new_Sorter100|18662_ ;
  assign \new_Sorter100|18763_  = \new_Sorter100|18663_  & \new_Sorter100|18664_ ;
  assign \new_Sorter100|18764_  = \new_Sorter100|18663_  | \new_Sorter100|18664_ ;
  assign \new_Sorter100|18765_  = \new_Sorter100|18665_  & \new_Sorter100|18666_ ;
  assign \new_Sorter100|18766_  = \new_Sorter100|18665_  | \new_Sorter100|18666_ ;
  assign \new_Sorter100|18767_  = \new_Sorter100|18667_  & \new_Sorter100|18668_ ;
  assign \new_Sorter100|18768_  = \new_Sorter100|18667_  | \new_Sorter100|18668_ ;
  assign \new_Sorter100|18769_  = \new_Sorter100|18669_  & \new_Sorter100|18670_ ;
  assign \new_Sorter100|18770_  = \new_Sorter100|18669_  | \new_Sorter100|18670_ ;
  assign \new_Sorter100|18771_  = \new_Sorter100|18671_  & \new_Sorter100|18672_ ;
  assign \new_Sorter100|18772_  = \new_Sorter100|18671_  | \new_Sorter100|18672_ ;
  assign \new_Sorter100|18773_  = \new_Sorter100|18673_  & \new_Sorter100|18674_ ;
  assign \new_Sorter100|18774_  = \new_Sorter100|18673_  | \new_Sorter100|18674_ ;
  assign \new_Sorter100|18775_  = \new_Sorter100|18675_  & \new_Sorter100|18676_ ;
  assign \new_Sorter100|18776_  = \new_Sorter100|18675_  | \new_Sorter100|18676_ ;
  assign \new_Sorter100|18777_  = \new_Sorter100|18677_  & \new_Sorter100|18678_ ;
  assign \new_Sorter100|18778_  = \new_Sorter100|18677_  | \new_Sorter100|18678_ ;
  assign \new_Sorter100|18779_  = \new_Sorter100|18679_  & \new_Sorter100|18680_ ;
  assign \new_Sorter100|18780_  = \new_Sorter100|18679_  | \new_Sorter100|18680_ ;
  assign \new_Sorter100|18781_  = \new_Sorter100|18681_  & \new_Sorter100|18682_ ;
  assign \new_Sorter100|18782_  = \new_Sorter100|18681_  | \new_Sorter100|18682_ ;
  assign \new_Sorter100|18783_  = \new_Sorter100|18683_  & \new_Sorter100|18684_ ;
  assign \new_Sorter100|18784_  = \new_Sorter100|18683_  | \new_Sorter100|18684_ ;
  assign \new_Sorter100|18785_  = \new_Sorter100|18685_  & \new_Sorter100|18686_ ;
  assign \new_Sorter100|18786_  = \new_Sorter100|18685_  | \new_Sorter100|18686_ ;
  assign \new_Sorter100|18787_  = \new_Sorter100|18687_  & \new_Sorter100|18688_ ;
  assign \new_Sorter100|18788_  = \new_Sorter100|18687_  | \new_Sorter100|18688_ ;
  assign \new_Sorter100|18789_  = \new_Sorter100|18689_  & \new_Sorter100|18690_ ;
  assign \new_Sorter100|18790_  = \new_Sorter100|18689_  | \new_Sorter100|18690_ ;
  assign \new_Sorter100|18791_  = \new_Sorter100|18691_  & \new_Sorter100|18692_ ;
  assign \new_Sorter100|18792_  = \new_Sorter100|18691_  | \new_Sorter100|18692_ ;
  assign \new_Sorter100|18793_  = \new_Sorter100|18693_  & \new_Sorter100|18694_ ;
  assign \new_Sorter100|18794_  = \new_Sorter100|18693_  | \new_Sorter100|18694_ ;
  assign \new_Sorter100|18795_  = \new_Sorter100|18695_  & \new_Sorter100|18696_ ;
  assign \new_Sorter100|18796_  = \new_Sorter100|18695_  | \new_Sorter100|18696_ ;
  assign \new_Sorter100|18797_  = \new_Sorter100|18697_  & \new_Sorter100|18698_ ;
  assign \new_Sorter100|18798_  = \new_Sorter100|18697_  | \new_Sorter100|18698_ ;
  assign \new_Sorter100|18800_  = \new_Sorter100|18700_  & \new_Sorter100|18701_ ;
  assign \new_Sorter100|18801_  = \new_Sorter100|18700_  | \new_Sorter100|18701_ ;
  assign \new_Sorter100|18802_  = \new_Sorter100|18702_  & \new_Sorter100|18703_ ;
  assign \new_Sorter100|18803_  = \new_Sorter100|18702_  | \new_Sorter100|18703_ ;
  assign \new_Sorter100|18804_  = \new_Sorter100|18704_  & \new_Sorter100|18705_ ;
  assign \new_Sorter100|18805_  = \new_Sorter100|18704_  | \new_Sorter100|18705_ ;
  assign \new_Sorter100|18806_  = \new_Sorter100|18706_  & \new_Sorter100|18707_ ;
  assign \new_Sorter100|18807_  = \new_Sorter100|18706_  | \new_Sorter100|18707_ ;
  assign \new_Sorter100|18808_  = \new_Sorter100|18708_  & \new_Sorter100|18709_ ;
  assign \new_Sorter100|18809_  = \new_Sorter100|18708_  | \new_Sorter100|18709_ ;
  assign \new_Sorter100|18810_  = \new_Sorter100|18710_  & \new_Sorter100|18711_ ;
  assign \new_Sorter100|18811_  = \new_Sorter100|18710_  | \new_Sorter100|18711_ ;
  assign \new_Sorter100|18812_  = \new_Sorter100|18712_  & \new_Sorter100|18713_ ;
  assign \new_Sorter100|18813_  = \new_Sorter100|18712_  | \new_Sorter100|18713_ ;
  assign \new_Sorter100|18814_  = \new_Sorter100|18714_  & \new_Sorter100|18715_ ;
  assign \new_Sorter100|18815_  = \new_Sorter100|18714_  | \new_Sorter100|18715_ ;
  assign \new_Sorter100|18816_  = \new_Sorter100|18716_  & \new_Sorter100|18717_ ;
  assign \new_Sorter100|18817_  = \new_Sorter100|18716_  | \new_Sorter100|18717_ ;
  assign \new_Sorter100|18818_  = \new_Sorter100|18718_  & \new_Sorter100|18719_ ;
  assign \new_Sorter100|18819_  = \new_Sorter100|18718_  | \new_Sorter100|18719_ ;
  assign \new_Sorter100|18820_  = \new_Sorter100|18720_  & \new_Sorter100|18721_ ;
  assign \new_Sorter100|18821_  = \new_Sorter100|18720_  | \new_Sorter100|18721_ ;
  assign \new_Sorter100|18822_  = \new_Sorter100|18722_  & \new_Sorter100|18723_ ;
  assign \new_Sorter100|18823_  = \new_Sorter100|18722_  | \new_Sorter100|18723_ ;
  assign \new_Sorter100|18824_  = \new_Sorter100|18724_  & \new_Sorter100|18725_ ;
  assign \new_Sorter100|18825_  = \new_Sorter100|18724_  | \new_Sorter100|18725_ ;
  assign \new_Sorter100|18826_  = \new_Sorter100|18726_  & \new_Sorter100|18727_ ;
  assign \new_Sorter100|18827_  = \new_Sorter100|18726_  | \new_Sorter100|18727_ ;
  assign \new_Sorter100|18828_  = \new_Sorter100|18728_  & \new_Sorter100|18729_ ;
  assign \new_Sorter100|18829_  = \new_Sorter100|18728_  | \new_Sorter100|18729_ ;
  assign \new_Sorter100|18830_  = \new_Sorter100|18730_  & \new_Sorter100|18731_ ;
  assign \new_Sorter100|18831_  = \new_Sorter100|18730_  | \new_Sorter100|18731_ ;
  assign \new_Sorter100|18832_  = \new_Sorter100|18732_  & \new_Sorter100|18733_ ;
  assign \new_Sorter100|18833_  = \new_Sorter100|18732_  | \new_Sorter100|18733_ ;
  assign \new_Sorter100|18834_  = \new_Sorter100|18734_  & \new_Sorter100|18735_ ;
  assign \new_Sorter100|18835_  = \new_Sorter100|18734_  | \new_Sorter100|18735_ ;
  assign \new_Sorter100|18836_  = \new_Sorter100|18736_  & \new_Sorter100|18737_ ;
  assign \new_Sorter100|18837_  = \new_Sorter100|18736_  | \new_Sorter100|18737_ ;
  assign \new_Sorter100|18838_  = \new_Sorter100|18738_  & \new_Sorter100|18739_ ;
  assign \new_Sorter100|18839_  = \new_Sorter100|18738_  | \new_Sorter100|18739_ ;
  assign \new_Sorter100|18840_  = \new_Sorter100|18740_  & \new_Sorter100|18741_ ;
  assign \new_Sorter100|18841_  = \new_Sorter100|18740_  | \new_Sorter100|18741_ ;
  assign \new_Sorter100|18842_  = \new_Sorter100|18742_  & \new_Sorter100|18743_ ;
  assign \new_Sorter100|18843_  = \new_Sorter100|18742_  | \new_Sorter100|18743_ ;
  assign \new_Sorter100|18844_  = \new_Sorter100|18744_  & \new_Sorter100|18745_ ;
  assign \new_Sorter100|18845_  = \new_Sorter100|18744_  | \new_Sorter100|18745_ ;
  assign \new_Sorter100|18846_  = \new_Sorter100|18746_  & \new_Sorter100|18747_ ;
  assign \new_Sorter100|18847_  = \new_Sorter100|18746_  | \new_Sorter100|18747_ ;
  assign \new_Sorter100|18848_  = \new_Sorter100|18748_  & \new_Sorter100|18749_ ;
  assign \new_Sorter100|18849_  = \new_Sorter100|18748_  | \new_Sorter100|18749_ ;
  assign \new_Sorter100|18850_  = \new_Sorter100|18750_  & \new_Sorter100|18751_ ;
  assign \new_Sorter100|18851_  = \new_Sorter100|18750_  | \new_Sorter100|18751_ ;
  assign \new_Sorter100|18852_  = \new_Sorter100|18752_  & \new_Sorter100|18753_ ;
  assign \new_Sorter100|18853_  = \new_Sorter100|18752_  | \new_Sorter100|18753_ ;
  assign \new_Sorter100|18854_  = \new_Sorter100|18754_  & \new_Sorter100|18755_ ;
  assign \new_Sorter100|18855_  = \new_Sorter100|18754_  | \new_Sorter100|18755_ ;
  assign \new_Sorter100|18856_  = \new_Sorter100|18756_  & \new_Sorter100|18757_ ;
  assign \new_Sorter100|18857_  = \new_Sorter100|18756_  | \new_Sorter100|18757_ ;
  assign \new_Sorter100|18858_  = \new_Sorter100|18758_  & \new_Sorter100|18759_ ;
  assign \new_Sorter100|18859_  = \new_Sorter100|18758_  | \new_Sorter100|18759_ ;
  assign \new_Sorter100|18860_  = \new_Sorter100|18760_  & \new_Sorter100|18761_ ;
  assign \new_Sorter100|18861_  = \new_Sorter100|18760_  | \new_Sorter100|18761_ ;
  assign \new_Sorter100|18862_  = \new_Sorter100|18762_  & \new_Sorter100|18763_ ;
  assign \new_Sorter100|18863_  = \new_Sorter100|18762_  | \new_Sorter100|18763_ ;
  assign \new_Sorter100|18864_  = \new_Sorter100|18764_  & \new_Sorter100|18765_ ;
  assign \new_Sorter100|18865_  = \new_Sorter100|18764_  | \new_Sorter100|18765_ ;
  assign \new_Sorter100|18866_  = \new_Sorter100|18766_  & \new_Sorter100|18767_ ;
  assign \new_Sorter100|18867_  = \new_Sorter100|18766_  | \new_Sorter100|18767_ ;
  assign \new_Sorter100|18868_  = \new_Sorter100|18768_  & \new_Sorter100|18769_ ;
  assign \new_Sorter100|18869_  = \new_Sorter100|18768_  | \new_Sorter100|18769_ ;
  assign \new_Sorter100|18870_  = \new_Sorter100|18770_  & \new_Sorter100|18771_ ;
  assign \new_Sorter100|18871_  = \new_Sorter100|18770_  | \new_Sorter100|18771_ ;
  assign \new_Sorter100|18872_  = \new_Sorter100|18772_  & \new_Sorter100|18773_ ;
  assign \new_Sorter100|18873_  = \new_Sorter100|18772_  | \new_Sorter100|18773_ ;
  assign \new_Sorter100|18874_  = \new_Sorter100|18774_  & \new_Sorter100|18775_ ;
  assign \new_Sorter100|18875_  = \new_Sorter100|18774_  | \new_Sorter100|18775_ ;
  assign \new_Sorter100|18876_  = \new_Sorter100|18776_  & \new_Sorter100|18777_ ;
  assign \new_Sorter100|18877_  = \new_Sorter100|18776_  | \new_Sorter100|18777_ ;
  assign \new_Sorter100|18878_  = \new_Sorter100|18778_  & \new_Sorter100|18779_ ;
  assign \new_Sorter100|18879_  = \new_Sorter100|18778_  | \new_Sorter100|18779_ ;
  assign \new_Sorter100|18880_  = \new_Sorter100|18780_  & \new_Sorter100|18781_ ;
  assign \new_Sorter100|18881_  = \new_Sorter100|18780_  | \new_Sorter100|18781_ ;
  assign \new_Sorter100|18882_  = \new_Sorter100|18782_  & \new_Sorter100|18783_ ;
  assign \new_Sorter100|18883_  = \new_Sorter100|18782_  | \new_Sorter100|18783_ ;
  assign \new_Sorter100|18884_  = \new_Sorter100|18784_  & \new_Sorter100|18785_ ;
  assign \new_Sorter100|18885_  = \new_Sorter100|18784_  | \new_Sorter100|18785_ ;
  assign \new_Sorter100|18886_  = \new_Sorter100|18786_  & \new_Sorter100|18787_ ;
  assign \new_Sorter100|18887_  = \new_Sorter100|18786_  | \new_Sorter100|18787_ ;
  assign \new_Sorter100|18888_  = \new_Sorter100|18788_  & \new_Sorter100|18789_ ;
  assign \new_Sorter100|18889_  = \new_Sorter100|18788_  | \new_Sorter100|18789_ ;
  assign \new_Sorter100|18890_  = \new_Sorter100|18790_  & \new_Sorter100|18791_ ;
  assign \new_Sorter100|18891_  = \new_Sorter100|18790_  | \new_Sorter100|18791_ ;
  assign \new_Sorter100|18892_  = \new_Sorter100|18792_  & \new_Sorter100|18793_ ;
  assign \new_Sorter100|18893_  = \new_Sorter100|18792_  | \new_Sorter100|18793_ ;
  assign \new_Sorter100|18894_  = \new_Sorter100|18794_  & \new_Sorter100|18795_ ;
  assign \new_Sorter100|18895_  = \new_Sorter100|18794_  | \new_Sorter100|18795_ ;
  assign \new_Sorter100|18896_  = \new_Sorter100|18796_  & \new_Sorter100|18797_ ;
  assign \new_Sorter100|18897_  = \new_Sorter100|18796_  | \new_Sorter100|18797_ ;
  assign \new_Sorter100|18898_  = \new_Sorter100|18798_  & \new_Sorter100|18799_ ;
  assign \new_Sorter100|18899_  = \new_Sorter100|18798_  | \new_Sorter100|18799_ ;
  assign \new_Sorter100|18900_  = \new_Sorter100|18800_ ;
  assign \new_Sorter100|18999_  = \new_Sorter100|18899_ ;
  assign \new_Sorter100|18901_  = \new_Sorter100|18801_  & \new_Sorter100|18802_ ;
  assign \new_Sorter100|18902_  = \new_Sorter100|18801_  | \new_Sorter100|18802_ ;
  assign \new_Sorter100|18903_  = \new_Sorter100|18803_  & \new_Sorter100|18804_ ;
  assign \new_Sorter100|18904_  = \new_Sorter100|18803_  | \new_Sorter100|18804_ ;
  assign \new_Sorter100|18905_  = \new_Sorter100|18805_  & \new_Sorter100|18806_ ;
  assign \new_Sorter100|18906_  = \new_Sorter100|18805_  | \new_Sorter100|18806_ ;
  assign \new_Sorter100|18907_  = \new_Sorter100|18807_  & \new_Sorter100|18808_ ;
  assign \new_Sorter100|18908_  = \new_Sorter100|18807_  | \new_Sorter100|18808_ ;
  assign \new_Sorter100|18909_  = \new_Sorter100|18809_  & \new_Sorter100|18810_ ;
  assign \new_Sorter100|18910_  = \new_Sorter100|18809_  | \new_Sorter100|18810_ ;
  assign \new_Sorter100|18911_  = \new_Sorter100|18811_  & \new_Sorter100|18812_ ;
  assign \new_Sorter100|18912_  = \new_Sorter100|18811_  | \new_Sorter100|18812_ ;
  assign \new_Sorter100|18913_  = \new_Sorter100|18813_  & \new_Sorter100|18814_ ;
  assign \new_Sorter100|18914_  = \new_Sorter100|18813_  | \new_Sorter100|18814_ ;
  assign \new_Sorter100|18915_  = \new_Sorter100|18815_  & \new_Sorter100|18816_ ;
  assign \new_Sorter100|18916_  = \new_Sorter100|18815_  | \new_Sorter100|18816_ ;
  assign \new_Sorter100|18917_  = \new_Sorter100|18817_  & \new_Sorter100|18818_ ;
  assign \new_Sorter100|18918_  = \new_Sorter100|18817_  | \new_Sorter100|18818_ ;
  assign \new_Sorter100|18919_  = \new_Sorter100|18819_  & \new_Sorter100|18820_ ;
  assign \new_Sorter100|18920_  = \new_Sorter100|18819_  | \new_Sorter100|18820_ ;
  assign \new_Sorter100|18921_  = \new_Sorter100|18821_  & \new_Sorter100|18822_ ;
  assign \new_Sorter100|18922_  = \new_Sorter100|18821_  | \new_Sorter100|18822_ ;
  assign \new_Sorter100|18923_  = \new_Sorter100|18823_  & \new_Sorter100|18824_ ;
  assign \new_Sorter100|18924_  = \new_Sorter100|18823_  | \new_Sorter100|18824_ ;
  assign \new_Sorter100|18925_  = \new_Sorter100|18825_  & \new_Sorter100|18826_ ;
  assign \new_Sorter100|18926_  = \new_Sorter100|18825_  | \new_Sorter100|18826_ ;
  assign \new_Sorter100|18927_  = \new_Sorter100|18827_  & \new_Sorter100|18828_ ;
  assign \new_Sorter100|18928_  = \new_Sorter100|18827_  | \new_Sorter100|18828_ ;
  assign \new_Sorter100|18929_  = \new_Sorter100|18829_  & \new_Sorter100|18830_ ;
  assign \new_Sorter100|18930_  = \new_Sorter100|18829_  | \new_Sorter100|18830_ ;
  assign \new_Sorter100|18931_  = \new_Sorter100|18831_  & \new_Sorter100|18832_ ;
  assign \new_Sorter100|18932_  = \new_Sorter100|18831_  | \new_Sorter100|18832_ ;
  assign \new_Sorter100|18933_  = \new_Sorter100|18833_  & \new_Sorter100|18834_ ;
  assign \new_Sorter100|18934_  = \new_Sorter100|18833_  | \new_Sorter100|18834_ ;
  assign \new_Sorter100|18935_  = \new_Sorter100|18835_  & \new_Sorter100|18836_ ;
  assign \new_Sorter100|18936_  = \new_Sorter100|18835_  | \new_Sorter100|18836_ ;
  assign \new_Sorter100|18937_  = \new_Sorter100|18837_  & \new_Sorter100|18838_ ;
  assign \new_Sorter100|18938_  = \new_Sorter100|18837_  | \new_Sorter100|18838_ ;
  assign \new_Sorter100|18939_  = \new_Sorter100|18839_  & \new_Sorter100|18840_ ;
  assign \new_Sorter100|18940_  = \new_Sorter100|18839_  | \new_Sorter100|18840_ ;
  assign \new_Sorter100|18941_  = \new_Sorter100|18841_  & \new_Sorter100|18842_ ;
  assign \new_Sorter100|18942_  = \new_Sorter100|18841_  | \new_Sorter100|18842_ ;
  assign \new_Sorter100|18943_  = \new_Sorter100|18843_  & \new_Sorter100|18844_ ;
  assign \new_Sorter100|18944_  = \new_Sorter100|18843_  | \new_Sorter100|18844_ ;
  assign \new_Sorter100|18945_  = \new_Sorter100|18845_  & \new_Sorter100|18846_ ;
  assign \new_Sorter100|18946_  = \new_Sorter100|18845_  | \new_Sorter100|18846_ ;
  assign \new_Sorter100|18947_  = \new_Sorter100|18847_  & \new_Sorter100|18848_ ;
  assign \new_Sorter100|18948_  = \new_Sorter100|18847_  | \new_Sorter100|18848_ ;
  assign \new_Sorter100|18949_  = \new_Sorter100|18849_  & \new_Sorter100|18850_ ;
  assign \new_Sorter100|18950_  = \new_Sorter100|18849_  | \new_Sorter100|18850_ ;
  assign \new_Sorter100|18951_  = \new_Sorter100|18851_  & \new_Sorter100|18852_ ;
  assign \new_Sorter100|18952_  = \new_Sorter100|18851_  | \new_Sorter100|18852_ ;
  assign \new_Sorter100|18953_  = \new_Sorter100|18853_  & \new_Sorter100|18854_ ;
  assign \new_Sorter100|18954_  = \new_Sorter100|18853_  | \new_Sorter100|18854_ ;
  assign \new_Sorter100|18955_  = \new_Sorter100|18855_  & \new_Sorter100|18856_ ;
  assign \new_Sorter100|18956_  = \new_Sorter100|18855_  | \new_Sorter100|18856_ ;
  assign \new_Sorter100|18957_  = \new_Sorter100|18857_  & \new_Sorter100|18858_ ;
  assign \new_Sorter100|18958_  = \new_Sorter100|18857_  | \new_Sorter100|18858_ ;
  assign \new_Sorter100|18959_  = \new_Sorter100|18859_  & \new_Sorter100|18860_ ;
  assign \new_Sorter100|18960_  = \new_Sorter100|18859_  | \new_Sorter100|18860_ ;
  assign \new_Sorter100|18961_  = \new_Sorter100|18861_  & \new_Sorter100|18862_ ;
  assign \new_Sorter100|18962_  = \new_Sorter100|18861_  | \new_Sorter100|18862_ ;
  assign \new_Sorter100|18963_  = \new_Sorter100|18863_  & \new_Sorter100|18864_ ;
  assign \new_Sorter100|18964_  = \new_Sorter100|18863_  | \new_Sorter100|18864_ ;
  assign \new_Sorter100|18965_  = \new_Sorter100|18865_  & \new_Sorter100|18866_ ;
  assign \new_Sorter100|18966_  = \new_Sorter100|18865_  | \new_Sorter100|18866_ ;
  assign \new_Sorter100|18967_  = \new_Sorter100|18867_  & \new_Sorter100|18868_ ;
  assign \new_Sorter100|18968_  = \new_Sorter100|18867_  | \new_Sorter100|18868_ ;
  assign \new_Sorter100|18969_  = \new_Sorter100|18869_  & \new_Sorter100|18870_ ;
  assign \new_Sorter100|18970_  = \new_Sorter100|18869_  | \new_Sorter100|18870_ ;
  assign \new_Sorter100|18971_  = \new_Sorter100|18871_  & \new_Sorter100|18872_ ;
  assign \new_Sorter100|18972_  = \new_Sorter100|18871_  | \new_Sorter100|18872_ ;
  assign \new_Sorter100|18973_  = \new_Sorter100|18873_  & \new_Sorter100|18874_ ;
  assign \new_Sorter100|18974_  = \new_Sorter100|18873_  | \new_Sorter100|18874_ ;
  assign \new_Sorter100|18975_  = \new_Sorter100|18875_  & \new_Sorter100|18876_ ;
  assign \new_Sorter100|18976_  = \new_Sorter100|18875_  | \new_Sorter100|18876_ ;
  assign \new_Sorter100|18977_  = \new_Sorter100|18877_  & \new_Sorter100|18878_ ;
  assign \new_Sorter100|18978_  = \new_Sorter100|18877_  | \new_Sorter100|18878_ ;
  assign \new_Sorter100|18979_  = \new_Sorter100|18879_  & \new_Sorter100|18880_ ;
  assign \new_Sorter100|18980_  = \new_Sorter100|18879_  | \new_Sorter100|18880_ ;
  assign \new_Sorter100|18981_  = \new_Sorter100|18881_  & \new_Sorter100|18882_ ;
  assign \new_Sorter100|18982_  = \new_Sorter100|18881_  | \new_Sorter100|18882_ ;
  assign \new_Sorter100|18983_  = \new_Sorter100|18883_  & \new_Sorter100|18884_ ;
  assign \new_Sorter100|18984_  = \new_Sorter100|18883_  | \new_Sorter100|18884_ ;
  assign \new_Sorter100|18985_  = \new_Sorter100|18885_  & \new_Sorter100|18886_ ;
  assign \new_Sorter100|18986_  = \new_Sorter100|18885_  | \new_Sorter100|18886_ ;
  assign \new_Sorter100|18987_  = \new_Sorter100|18887_  & \new_Sorter100|18888_ ;
  assign \new_Sorter100|18988_  = \new_Sorter100|18887_  | \new_Sorter100|18888_ ;
  assign \new_Sorter100|18989_  = \new_Sorter100|18889_  & \new_Sorter100|18890_ ;
  assign \new_Sorter100|18990_  = \new_Sorter100|18889_  | \new_Sorter100|18890_ ;
  assign \new_Sorter100|18991_  = \new_Sorter100|18891_  & \new_Sorter100|18892_ ;
  assign \new_Sorter100|18992_  = \new_Sorter100|18891_  | \new_Sorter100|18892_ ;
  assign \new_Sorter100|18993_  = \new_Sorter100|18893_  & \new_Sorter100|18894_ ;
  assign \new_Sorter100|18994_  = \new_Sorter100|18893_  | \new_Sorter100|18894_ ;
  assign \new_Sorter100|18995_  = \new_Sorter100|18895_  & \new_Sorter100|18896_ ;
  assign \new_Sorter100|18996_  = \new_Sorter100|18895_  | \new_Sorter100|18896_ ;
  assign \new_Sorter100|18997_  = \new_Sorter100|18897_  & \new_Sorter100|18898_ ;
  assign \new_Sorter100|18998_  = \new_Sorter100|18897_  | \new_Sorter100|18898_ ;
  assign \new_Sorter100|19000_  = \new_Sorter100|18900_  & \new_Sorter100|18901_ ;
  assign \new_Sorter100|19001_  = \new_Sorter100|18900_  | \new_Sorter100|18901_ ;
  assign \new_Sorter100|19002_  = \new_Sorter100|18902_  & \new_Sorter100|18903_ ;
  assign \new_Sorter100|19003_  = \new_Sorter100|18902_  | \new_Sorter100|18903_ ;
  assign \new_Sorter100|19004_  = \new_Sorter100|18904_  & \new_Sorter100|18905_ ;
  assign \new_Sorter100|19005_  = \new_Sorter100|18904_  | \new_Sorter100|18905_ ;
  assign \new_Sorter100|19006_  = \new_Sorter100|18906_  & \new_Sorter100|18907_ ;
  assign \new_Sorter100|19007_  = \new_Sorter100|18906_  | \new_Sorter100|18907_ ;
  assign \new_Sorter100|19008_  = \new_Sorter100|18908_  & \new_Sorter100|18909_ ;
  assign \new_Sorter100|19009_  = \new_Sorter100|18908_  | \new_Sorter100|18909_ ;
  assign \new_Sorter100|19010_  = \new_Sorter100|18910_  & \new_Sorter100|18911_ ;
  assign \new_Sorter100|19011_  = \new_Sorter100|18910_  | \new_Sorter100|18911_ ;
  assign \new_Sorter100|19012_  = \new_Sorter100|18912_  & \new_Sorter100|18913_ ;
  assign \new_Sorter100|19013_  = \new_Sorter100|18912_  | \new_Sorter100|18913_ ;
  assign \new_Sorter100|19014_  = \new_Sorter100|18914_  & \new_Sorter100|18915_ ;
  assign \new_Sorter100|19015_  = \new_Sorter100|18914_  | \new_Sorter100|18915_ ;
  assign \new_Sorter100|19016_  = \new_Sorter100|18916_  & \new_Sorter100|18917_ ;
  assign \new_Sorter100|19017_  = \new_Sorter100|18916_  | \new_Sorter100|18917_ ;
  assign \new_Sorter100|19018_  = \new_Sorter100|18918_  & \new_Sorter100|18919_ ;
  assign \new_Sorter100|19019_  = \new_Sorter100|18918_  | \new_Sorter100|18919_ ;
  assign \new_Sorter100|19020_  = \new_Sorter100|18920_  & \new_Sorter100|18921_ ;
  assign \new_Sorter100|19021_  = \new_Sorter100|18920_  | \new_Sorter100|18921_ ;
  assign \new_Sorter100|19022_  = \new_Sorter100|18922_  & \new_Sorter100|18923_ ;
  assign \new_Sorter100|19023_  = \new_Sorter100|18922_  | \new_Sorter100|18923_ ;
  assign \new_Sorter100|19024_  = \new_Sorter100|18924_  & \new_Sorter100|18925_ ;
  assign \new_Sorter100|19025_  = \new_Sorter100|18924_  | \new_Sorter100|18925_ ;
  assign \new_Sorter100|19026_  = \new_Sorter100|18926_  & \new_Sorter100|18927_ ;
  assign \new_Sorter100|19027_  = \new_Sorter100|18926_  | \new_Sorter100|18927_ ;
  assign \new_Sorter100|19028_  = \new_Sorter100|18928_  & \new_Sorter100|18929_ ;
  assign \new_Sorter100|19029_  = \new_Sorter100|18928_  | \new_Sorter100|18929_ ;
  assign \new_Sorter100|19030_  = \new_Sorter100|18930_  & \new_Sorter100|18931_ ;
  assign \new_Sorter100|19031_  = \new_Sorter100|18930_  | \new_Sorter100|18931_ ;
  assign \new_Sorter100|19032_  = \new_Sorter100|18932_  & \new_Sorter100|18933_ ;
  assign \new_Sorter100|19033_  = \new_Sorter100|18932_  | \new_Sorter100|18933_ ;
  assign \new_Sorter100|19034_  = \new_Sorter100|18934_  & \new_Sorter100|18935_ ;
  assign \new_Sorter100|19035_  = \new_Sorter100|18934_  | \new_Sorter100|18935_ ;
  assign \new_Sorter100|19036_  = \new_Sorter100|18936_  & \new_Sorter100|18937_ ;
  assign \new_Sorter100|19037_  = \new_Sorter100|18936_  | \new_Sorter100|18937_ ;
  assign \new_Sorter100|19038_  = \new_Sorter100|18938_  & \new_Sorter100|18939_ ;
  assign \new_Sorter100|19039_  = \new_Sorter100|18938_  | \new_Sorter100|18939_ ;
  assign \new_Sorter100|19040_  = \new_Sorter100|18940_  & \new_Sorter100|18941_ ;
  assign \new_Sorter100|19041_  = \new_Sorter100|18940_  | \new_Sorter100|18941_ ;
  assign \new_Sorter100|19042_  = \new_Sorter100|18942_  & \new_Sorter100|18943_ ;
  assign \new_Sorter100|19043_  = \new_Sorter100|18942_  | \new_Sorter100|18943_ ;
  assign \new_Sorter100|19044_  = \new_Sorter100|18944_  & \new_Sorter100|18945_ ;
  assign \new_Sorter100|19045_  = \new_Sorter100|18944_  | \new_Sorter100|18945_ ;
  assign \new_Sorter100|19046_  = \new_Sorter100|18946_  & \new_Sorter100|18947_ ;
  assign \new_Sorter100|19047_  = \new_Sorter100|18946_  | \new_Sorter100|18947_ ;
  assign \new_Sorter100|19048_  = \new_Sorter100|18948_  & \new_Sorter100|18949_ ;
  assign \new_Sorter100|19049_  = \new_Sorter100|18948_  | \new_Sorter100|18949_ ;
  assign \new_Sorter100|19050_  = \new_Sorter100|18950_  & \new_Sorter100|18951_ ;
  assign \new_Sorter100|19051_  = \new_Sorter100|18950_  | \new_Sorter100|18951_ ;
  assign \new_Sorter100|19052_  = \new_Sorter100|18952_  & \new_Sorter100|18953_ ;
  assign \new_Sorter100|19053_  = \new_Sorter100|18952_  | \new_Sorter100|18953_ ;
  assign \new_Sorter100|19054_  = \new_Sorter100|18954_  & \new_Sorter100|18955_ ;
  assign \new_Sorter100|19055_  = \new_Sorter100|18954_  | \new_Sorter100|18955_ ;
  assign \new_Sorter100|19056_  = \new_Sorter100|18956_  & \new_Sorter100|18957_ ;
  assign \new_Sorter100|19057_  = \new_Sorter100|18956_  | \new_Sorter100|18957_ ;
  assign \new_Sorter100|19058_  = \new_Sorter100|18958_  & \new_Sorter100|18959_ ;
  assign \new_Sorter100|19059_  = \new_Sorter100|18958_  | \new_Sorter100|18959_ ;
  assign \new_Sorter100|19060_  = \new_Sorter100|18960_  & \new_Sorter100|18961_ ;
  assign \new_Sorter100|19061_  = \new_Sorter100|18960_  | \new_Sorter100|18961_ ;
  assign \new_Sorter100|19062_  = \new_Sorter100|18962_  & \new_Sorter100|18963_ ;
  assign \new_Sorter100|19063_  = \new_Sorter100|18962_  | \new_Sorter100|18963_ ;
  assign \new_Sorter100|19064_  = \new_Sorter100|18964_  & \new_Sorter100|18965_ ;
  assign \new_Sorter100|19065_  = \new_Sorter100|18964_  | \new_Sorter100|18965_ ;
  assign \new_Sorter100|19066_  = \new_Sorter100|18966_  & \new_Sorter100|18967_ ;
  assign \new_Sorter100|19067_  = \new_Sorter100|18966_  | \new_Sorter100|18967_ ;
  assign \new_Sorter100|19068_  = \new_Sorter100|18968_  & \new_Sorter100|18969_ ;
  assign \new_Sorter100|19069_  = \new_Sorter100|18968_  | \new_Sorter100|18969_ ;
  assign \new_Sorter100|19070_  = \new_Sorter100|18970_  & \new_Sorter100|18971_ ;
  assign \new_Sorter100|19071_  = \new_Sorter100|18970_  | \new_Sorter100|18971_ ;
  assign \new_Sorter100|19072_  = \new_Sorter100|18972_  & \new_Sorter100|18973_ ;
  assign \new_Sorter100|19073_  = \new_Sorter100|18972_  | \new_Sorter100|18973_ ;
  assign \new_Sorter100|19074_  = \new_Sorter100|18974_  & \new_Sorter100|18975_ ;
  assign \new_Sorter100|19075_  = \new_Sorter100|18974_  | \new_Sorter100|18975_ ;
  assign \new_Sorter100|19076_  = \new_Sorter100|18976_  & \new_Sorter100|18977_ ;
  assign \new_Sorter100|19077_  = \new_Sorter100|18976_  | \new_Sorter100|18977_ ;
  assign \new_Sorter100|19078_  = \new_Sorter100|18978_  & \new_Sorter100|18979_ ;
  assign \new_Sorter100|19079_  = \new_Sorter100|18978_  | \new_Sorter100|18979_ ;
  assign \new_Sorter100|19080_  = \new_Sorter100|18980_  & \new_Sorter100|18981_ ;
  assign \new_Sorter100|19081_  = \new_Sorter100|18980_  | \new_Sorter100|18981_ ;
  assign \new_Sorter100|19082_  = \new_Sorter100|18982_  & \new_Sorter100|18983_ ;
  assign \new_Sorter100|19083_  = \new_Sorter100|18982_  | \new_Sorter100|18983_ ;
  assign \new_Sorter100|19084_  = \new_Sorter100|18984_  & \new_Sorter100|18985_ ;
  assign \new_Sorter100|19085_  = \new_Sorter100|18984_  | \new_Sorter100|18985_ ;
  assign \new_Sorter100|19086_  = \new_Sorter100|18986_  & \new_Sorter100|18987_ ;
  assign \new_Sorter100|19087_  = \new_Sorter100|18986_  | \new_Sorter100|18987_ ;
  assign \new_Sorter100|19088_  = \new_Sorter100|18988_  & \new_Sorter100|18989_ ;
  assign \new_Sorter100|19089_  = \new_Sorter100|18988_  | \new_Sorter100|18989_ ;
  assign \new_Sorter100|19090_  = \new_Sorter100|18990_  & \new_Sorter100|18991_ ;
  assign \new_Sorter100|19091_  = \new_Sorter100|18990_  | \new_Sorter100|18991_ ;
  assign \new_Sorter100|19092_  = \new_Sorter100|18992_  & \new_Sorter100|18993_ ;
  assign \new_Sorter100|19093_  = \new_Sorter100|18992_  | \new_Sorter100|18993_ ;
  assign \new_Sorter100|19094_  = \new_Sorter100|18994_  & \new_Sorter100|18995_ ;
  assign \new_Sorter100|19095_  = \new_Sorter100|18994_  | \new_Sorter100|18995_ ;
  assign \new_Sorter100|19096_  = \new_Sorter100|18996_  & \new_Sorter100|18997_ ;
  assign \new_Sorter100|19097_  = \new_Sorter100|18996_  | \new_Sorter100|18997_ ;
  assign \new_Sorter100|19098_  = \new_Sorter100|18998_  & \new_Sorter100|18999_ ;
  assign \new_Sorter100|19099_  = \new_Sorter100|18998_  | \new_Sorter100|18999_ ;
  assign \new_Sorter100|19100_  = \new_Sorter100|19000_ ;
  assign \new_Sorter100|19199_  = \new_Sorter100|19099_ ;
  assign \new_Sorter100|19101_  = \new_Sorter100|19001_  & \new_Sorter100|19002_ ;
  assign \new_Sorter100|19102_  = \new_Sorter100|19001_  | \new_Sorter100|19002_ ;
  assign \new_Sorter100|19103_  = \new_Sorter100|19003_  & \new_Sorter100|19004_ ;
  assign \new_Sorter100|19104_  = \new_Sorter100|19003_  | \new_Sorter100|19004_ ;
  assign \new_Sorter100|19105_  = \new_Sorter100|19005_  & \new_Sorter100|19006_ ;
  assign \new_Sorter100|19106_  = \new_Sorter100|19005_  | \new_Sorter100|19006_ ;
  assign \new_Sorter100|19107_  = \new_Sorter100|19007_  & \new_Sorter100|19008_ ;
  assign \new_Sorter100|19108_  = \new_Sorter100|19007_  | \new_Sorter100|19008_ ;
  assign \new_Sorter100|19109_  = \new_Sorter100|19009_  & \new_Sorter100|19010_ ;
  assign \new_Sorter100|19110_  = \new_Sorter100|19009_  | \new_Sorter100|19010_ ;
  assign \new_Sorter100|19111_  = \new_Sorter100|19011_  & \new_Sorter100|19012_ ;
  assign \new_Sorter100|19112_  = \new_Sorter100|19011_  | \new_Sorter100|19012_ ;
  assign \new_Sorter100|19113_  = \new_Sorter100|19013_  & \new_Sorter100|19014_ ;
  assign \new_Sorter100|19114_  = \new_Sorter100|19013_  | \new_Sorter100|19014_ ;
  assign \new_Sorter100|19115_  = \new_Sorter100|19015_  & \new_Sorter100|19016_ ;
  assign \new_Sorter100|19116_  = \new_Sorter100|19015_  | \new_Sorter100|19016_ ;
  assign \new_Sorter100|19117_  = \new_Sorter100|19017_  & \new_Sorter100|19018_ ;
  assign \new_Sorter100|19118_  = \new_Sorter100|19017_  | \new_Sorter100|19018_ ;
  assign \new_Sorter100|19119_  = \new_Sorter100|19019_  & \new_Sorter100|19020_ ;
  assign \new_Sorter100|19120_  = \new_Sorter100|19019_  | \new_Sorter100|19020_ ;
  assign \new_Sorter100|19121_  = \new_Sorter100|19021_  & \new_Sorter100|19022_ ;
  assign \new_Sorter100|19122_  = \new_Sorter100|19021_  | \new_Sorter100|19022_ ;
  assign \new_Sorter100|19123_  = \new_Sorter100|19023_  & \new_Sorter100|19024_ ;
  assign \new_Sorter100|19124_  = \new_Sorter100|19023_  | \new_Sorter100|19024_ ;
  assign \new_Sorter100|19125_  = \new_Sorter100|19025_  & \new_Sorter100|19026_ ;
  assign \new_Sorter100|19126_  = \new_Sorter100|19025_  | \new_Sorter100|19026_ ;
  assign \new_Sorter100|19127_  = \new_Sorter100|19027_  & \new_Sorter100|19028_ ;
  assign \new_Sorter100|19128_  = \new_Sorter100|19027_  | \new_Sorter100|19028_ ;
  assign \new_Sorter100|19129_  = \new_Sorter100|19029_  & \new_Sorter100|19030_ ;
  assign \new_Sorter100|19130_  = \new_Sorter100|19029_  | \new_Sorter100|19030_ ;
  assign \new_Sorter100|19131_  = \new_Sorter100|19031_  & \new_Sorter100|19032_ ;
  assign \new_Sorter100|19132_  = \new_Sorter100|19031_  | \new_Sorter100|19032_ ;
  assign \new_Sorter100|19133_  = \new_Sorter100|19033_  & \new_Sorter100|19034_ ;
  assign \new_Sorter100|19134_  = \new_Sorter100|19033_  | \new_Sorter100|19034_ ;
  assign \new_Sorter100|19135_  = \new_Sorter100|19035_  & \new_Sorter100|19036_ ;
  assign \new_Sorter100|19136_  = \new_Sorter100|19035_  | \new_Sorter100|19036_ ;
  assign \new_Sorter100|19137_  = \new_Sorter100|19037_  & \new_Sorter100|19038_ ;
  assign \new_Sorter100|19138_  = \new_Sorter100|19037_  | \new_Sorter100|19038_ ;
  assign \new_Sorter100|19139_  = \new_Sorter100|19039_  & \new_Sorter100|19040_ ;
  assign \new_Sorter100|19140_  = \new_Sorter100|19039_  | \new_Sorter100|19040_ ;
  assign \new_Sorter100|19141_  = \new_Sorter100|19041_  & \new_Sorter100|19042_ ;
  assign \new_Sorter100|19142_  = \new_Sorter100|19041_  | \new_Sorter100|19042_ ;
  assign \new_Sorter100|19143_  = \new_Sorter100|19043_  & \new_Sorter100|19044_ ;
  assign \new_Sorter100|19144_  = \new_Sorter100|19043_  | \new_Sorter100|19044_ ;
  assign \new_Sorter100|19145_  = \new_Sorter100|19045_  & \new_Sorter100|19046_ ;
  assign \new_Sorter100|19146_  = \new_Sorter100|19045_  | \new_Sorter100|19046_ ;
  assign \new_Sorter100|19147_  = \new_Sorter100|19047_  & \new_Sorter100|19048_ ;
  assign \new_Sorter100|19148_  = \new_Sorter100|19047_  | \new_Sorter100|19048_ ;
  assign \new_Sorter100|19149_  = \new_Sorter100|19049_  & \new_Sorter100|19050_ ;
  assign \new_Sorter100|19150_  = \new_Sorter100|19049_  | \new_Sorter100|19050_ ;
  assign \new_Sorter100|19151_  = \new_Sorter100|19051_  & \new_Sorter100|19052_ ;
  assign \new_Sorter100|19152_  = \new_Sorter100|19051_  | \new_Sorter100|19052_ ;
  assign \new_Sorter100|19153_  = \new_Sorter100|19053_  & \new_Sorter100|19054_ ;
  assign \new_Sorter100|19154_  = \new_Sorter100|19053_  | \new_Sorter100|19054_ ;
  assign \new_Sorter100|19155_  = \new_Sorter100|19055_  & \new_Sorter100|19056_ ;
  assign \new_Sorter100|19156_  = \new_Sorter100|19055_  | \new_Sorter100|19056_ ;
  assign \new_Sorter100|19157_  = \new_Sorter100|19057_  & \new_Sorter100|19058_ ;
  assign \new_Sorter100|19158_  = \new_Sorter100|19057_  | \new_Sorter100|19058_ ;
  assign \new_Sorter100|19159_  = \new_Sorter100|19059_  & \new_Sorter100|19060_ ;
  assign \new_Sorter100|19160_  = \new_Sorter100|19059_  | \new_Sorter100|19060_ ;
  assign \new_Sorter100|19161_  = \new_Sorter100|19061_  & \new_Sorter100|19062_ ;
  assign \new_Sorter100|19162_  = \new_Sorter100|19061_  | \new_Sorter100|19062_ ;
  assign \new_Sorter100|19163_  = \new_Sorter100|19063_  & \new_Sorter100|19064_ ;
  assign \new_Sorter100|19164_  = \new_Sorter100|19063_  | \new_Sorter100|19064_ ;
  assign \new_Sorter100|19165_  = \new_Sorter100|19065_  & \new_Sorter100|19066_ ;
  assign \new_Sorter100|19166_  = \new_Sorter100|19065_  | \new_Sorter100|19066_ ;
  assign \new_Sorter100|19167_  = \new_Sorter100|19067_  & \new_Sorter100|19068_ ;
  assign \new_Sorter100|19168_  = \new_Sorter100|19067_  | \new_Sorter100|19068_ ;
  assign \new_Sorter100|19169_  = \new_Sorter100|19069_  & \new_Sorter100|19070_ ;
  assign \new_Sorter100|19170_  = \new_Sorter100|19069_  | \new_Sorter100|19070_ ;
  assign \new_Sorter100|19171_  = \new_Sorter100|19071_  & \new_Sorter100|19072_ ;
  assign \new_Sorter100|19172_  = \new_Sorter100|19071_  | \new_Sorter100|19072_ ;
  assign \new_Sorter100|19173_  = \new_Sorter100|19073_  & \new_Sorter100|19074_ ;
  assign \new_Sorter100|19174_  = \new_Sorter100|19073_  | \new_Sorter100|19074_ ;
  assign \new_Sorter100|19175_  = \new_Sorter100|19075_  & \new_Sorter100|19076_ ;
  assign \new_Sorter100|19176_  = \new_Sorter100|19075_  | \new_Sorter100|19076_ ;
  assign \new_Sorter100|19177_  = \new_Sorter100|19077_  & \new_Sorter100|19078_ ;
  assign \new_Sorter100|19178_  = \new_Sorter100|19077_  | \new_Sorter100|19078_ ;
  assign \new_Sorter100|19179_  = \new_Sorter100|19079_  & \new_Sorter100|19080_ ;
  assign \new_Sorter100|19180_  = \new_Sorter100|19079_  | \new_Sorter100|19080_ ;
  assign \new_Sorter100|19181_  = \new_Sorter100|19081_  & \new_Sorter100|19082_ ;
  assign \new_Sorter100|19182_  = \new_Sorter100|19081_  | \new_Sorter100|19082_ ;
  assign \new_Sorter100|19183_  = \new_Sorter100|19083_  & \new_Sorter100|19084_ ;
  assign \new_Sorter100|19184_  = \new_Sorter100|19083_  | \new_Sorter100|19084_ ;
  assign \new_Sorter100|19185_  = \new_Sorter100|19085_  & \new_Sorter100|19086_ ;
  assign \new_Sorter100|19186_  = \new_Sorter100|19085_  | \new_Sorter100|19086_ ;
  assign \new_Sorter100|19187_  = \new_Sorter100|19087_  & \new_Sorter100|19088_ ;
  assign \new_Sorter100|19188_  = \new_Sorter100|19087_  | \new_Sorter100|19088_ ;
  assign \new_Sorter100|19189_  = \new_Sorter100|19089_  & \new_Sorter100|19090_ ;
  assign \new_Sorter100|19190_  = \new_Sorter100|19089_  | \new_Sorter100|19090_ ;
  assign \new_Sorter100|19191_  = \new_Sorter100|19091_  & \new_Sorter100|19092_ ;
  assign \new_Sorter100|19192_  = \new_Sorter100|19091_  | \new_Sorter100|19092_ ;
  assign \new_Sorter100|19193_  = \new_Sorter100|19093_  & \new_Sorter100|19094_ ;
  assign \new_Sorter100|19194_  = \new_Sorter100|19093_  | \new_Sorter100|19094_ ;
  assign \new_Sorter100|19195_  = \new_Sorter100|19095_  & \new_Sorter100|19096_ ;
  assign \new_Sorter100|19196_  = \new_Sorter100|19095_  | \new_Sorter100|19096_ ;
  assign \new_Sorter100|19197_  = \new_Sorter100|19097_  & \new_Sorter100|19098_ ;
  assign \new_Sorter100|19198_  = \new_Sorter100|19097_  | \new_Sorter100|19098_ ;
  assign \new_Sorter100|19200_  = \new_Sorter100|19100_  & \new_Sorter100|19101_ ;
  assign \new_Sorter100|19201_  = \new_Sorter100|19100_  | \new_Sorter100|19101_ ;
  assign \new_Sorter100|19202_  = \new_Sorter100|19102_  & \new_Sorter100|19103_ ;
  assign \new_Sorter100|19203_  = \new_Sorter100|19102_  | \new_Sorter100|19103_ ;
  assign \new_Sorter100|19204_  = \new_Sorter100|19104_  & \new_Sorter100|19105_ ;
  assign \new_Sorter100|19205_  = \new_Sorter100|19104_  | \new_Sorter100|19105_ ;
  assign \new_Sorter100|19206_  = \new_Sorter100|19106_  & \new_Sorter100|19107_ ;
  assign \new_Sorter100|19207_  = \new_Sorter100|19106_  | \new_Sorter100|19107_ ;
  assign \new_Sorter100|19208_  = \new_Sorter100|19108_  & \new_Sorter100|19109_ ;
  assign \new_Sorter100|19209_  = \new_Sorter100|19108_  | \new_Sorter100|19109_ ;
  assign \new_Sorter100|19210_  = \new_Sorter100|19110_  & \new_Sorter100|19111_ ;
  assign \new_Sorter100|19211_  = \new_Sorter100|19110_  | \new_Sorter100|19111_ ;
  assign \new_Sorter100|19212_  = \new_Sorter100|19112_  & \new_Sorter100|19113_ ;
  assign \new_Sorter100|19213_  = \new_Sorter100|19112_  | \new_Sorter100|19113_ ;
  assign \new_Sorter100|19214_  = \new_Sorter100|19114_  & \new_Sorter100|19115_ ;
  assign \new_Sorter100|19215_  = \new_Sorter100|19114_  | \new_Sorter100|19115_ ;
  assign \new_Sorter100|19216_  = \new_Sorter100|19116_  & \new_Sorter100|19117_ ;
  assign \new_Sorter100|19217_  = \new_Sorter100|19116_  | \new_Sorter100|19117_ ;
  assign \new_Sorter100|19218_  = \new_Sorter100|19118_  & \new_Sorter100|19119_ ;
  assign \new_Sorter100|19219_  = \new_Sorter100|19118_  | \new_Sorter100|19119_ ;
  assign \new_Sorter100|19220_  = \new_Sorter100|19120_  & \new_Sorter100|19121_ ;
  assign \new_Sorter100|19221_  = \new_Sorter100|19120_  | \new_Sorter100|19121_ ;
  assign \new_Sorter100|19222_  = \new_Sorter100|19122_  & \new_Sorter100|19123_ ;
  assign \new_Sorter100|19223_  = \new_Sorter100|19122_  | \new_Sorter100|19123_ ;
  assign \new_Sorter100|19224_  = \new_Sorter100|19124_  & \new_Sorter100|19125_ ;
  assign \new_Sorter100|19225_  = \new_Sorter100|19124_  | \new_Sorter100|19125_ ;
  assign \new_Sorter100|19226_  = \new_Sorter100|19126_  & \new_Sorter100|19127_ ;
  assign \new_Sorter100|19227_  = \new_Sorter100|19126_  | \new_Sorter100|19127_ ;
  assign \new_Sorter100|19228_  = \new_Sorter100|19128_  & \new_Sorter100|19129_ ;
  assign \new_Sorter100|19229_  = \new_Sorter100|19128_  | \new_Sorter100|19129_ ;
  assign \new_Sorter100|19230_  = \new_Sorter100|19130_  & \new_Sorter100|19131_ ;
  assign \new_Sorter100|19231_  = \new_Sorter100|19130_  | \new_Sorter100|19131_ ;
  assign \new_Sorter100|19232_  = \new_Sorter100|19132_  & \new_Sorter100|19133_ ;
  assign \new_Sorter100|19233_  = \new_Sorter100|19132_  | \new_Sorter100|19133_ ;
  assign \new_Sorter100|19234_  = \new_Sorter100|19134_  & \new_Sorter100|19135_ ;
  assign \new_Sorter100|19235_  = \new_Sorter100|19134_  | \new_Sorter100|19135_ ;
  assign \new_Sorter100|19236_  = \new_Sorter100|19136_  & \new_Sorter100|19137_ ;
  assign \new_Sorter100|19237_  = \new_Sorter100|19136_  | \new_Sorter100|19137_ ;
  assign \new_Sorter100|19238_  = \new_Sorter100|19138_  & \new_Sorter100|19139_ ;
  assign \new_Sorter100|19239_  = \new_Sorter100|19138_  | \new_Sorter100|19139_ ;
  assign \new_Sorter100|19240_  = \new_Sorter100|19140_  & \new_Sorter100|19141_ ;
  assign \new_Sorter100|19241_  = \new_Sorter100|19140_  | \new_Sorter100|19141_ ;
  assign \new_Sorter100|19242_  = \new_Sorter100|19142_  & \new_Sorter100|19143_ ;
  assign \new_Sorter100|19243_  = \new_Sorter100|19142_  | \new_Sorter100|19143_ ;
  assign \new_Sorter100|19244_  = \new_Sorter100|19144_  & \new_Sorter100|19145_ ;
  assign \new_Sorter100|19245_  = \new_Sorter100|19144_  | \new_Sorter100|19145_ ;
  assign \new_Sorter100|19246_  = \new_Sorter100|19146_  & \new_Sorter100|19147_ ;
  assign \new_Sorter100|19247_  = \new_Sorter100|19146_  | \new_Sorter100|19147_ ;
  assign \new_Sorter100|19248_  = \new_Sorter100|19148_  & \new_Sorter100|19149_ ;
  assign \new_Sorter100|19249_  = \new_Sorter100|19148_  | \new_Sorter100|19149_ ;
  assign \new_Sorter100|19250_  = \new_Sorter100|19150_  & \new_Sorter100|19151_ ;
  assign \new_Sorter100|19251_  = \new_Sorter100|19150_  | \new_Sorter100|19151_ ;
  assign \new_Sorter100|19252_  = \new_Sorter100|19152_  & \new_Sorter100|19153_ ;
  assign \new_Sorter100|19253_  = \new_Sorter100|19152_  | \new_Sorter100|19153_ ;
  assign \new_Sorter100|19254_  = \new_Sorter100|19154_  & \new_Sorter100|19155_ ;
  assign \new_Sorter100|19255_  = \new_Sorter100|19154_  | \new_Sorter100|19155_ ;
  assign \new_Sorter100|19256_  = \new_Sorter100|19156_  & \new_Sorter100|19157_ ;
  assign \new_Sorter100|19257_  = \new_Sorter100|19156_  | \new_Sorter100|19157_ ;
  assign \new_Sorter100|19258_  = \new_Sorter100|19158_  & \new_Sorter100|19159_ ;
  assign \new_Sorter100|19259_  = \new_Sorter100|19158_  | \new_Sorter100|19159_ ;
  assign \new_Sorter100|19260_  = \new_Sorter100|19160_  & \new_Sorter100|19161_ ;
  assign \new_Sorter100|19261_  = \new_Sorter100|19160_  | \new_Sorter100|19161_ ;
  assign \new_Sorter100|19262_  = \new_Sorter100|19162_  & \new_Sorter100|19163_ ;
  assign \new_Sorter100|19263_  = \new_Sorter100|19162_  | \new_Sorter100|19163_ ;
  assign \new_Sorter100|19264_  = \new_Sorter100|19164_  & \new_Sorter100|19165_ ;
  assign \new_Sorter100|19265_  = \new_Sorter100|19164_  | \new_Sorter100|19165_ ;
  assign \new_Sorter100|19266_  = \new_Sorter100|19166_  & \new_Sorter100|19167_ ;
  assign \new_Sorter100|19267_  = \new_Sorter100|19166_  | \new_Sorter100|19167_ ;
  assign \new_Sorter100|19268_  = \new_Sorter100|19168_  & \new_Sorter100|19169_ ;
  assign \new_Sorter100|19269_  = \new_Sorter100|19168_  | \new_Sorter100|19169_ ;
  assign \new_Sorter100|19270_  = \new_Sorter100|19170_  & \new_Sorter100|19171_ ;
  assign \new_Sorter100|19271_  = \new_Sorter100|19170_  | \new_Sorter100|19171_ ;
  assign \new_Sorter100|19272_  = \new_Sorter100|19172_  & \new_Sorter100|19173_ ;
  assign \new_Sorter100|19273_  = \new_Sorter100|19172_  | \new_Sorter100|19173_ ;
  assign \new_Sorter100|19274_  = \new_Sorter100|19174_  & \new_Sorter100|19175_ ;
  assign \new_Sorter100|19275_  = \new_Sorter100|19174_  | \new_Sorter100|19175_ ;
  assign \new_Sorter100|19276_  = \new_Sorter100|19176_  & \new_Sorter100|19177_ ;
  assign \new_Sorter100|19277_  = \new_Sorter100|19176_  | \new_Sorter100|19177_ ;
  assign \new_Sorter100|19278_  = \new_Sorter100|19178_  & \new_Sorter100|19179_ ;
  assign \new_Sorter100|19279_  = \new_Sorter100|19178_  | \new_Sorter100|19179_ ;
  assign \new_Sorter100|19280_  = \new_Sorter100|19180_  & \new_Sorter100|19181_ ;
  assign \new_Sorter100|19281_  = \new_Sorter100|19180_  | \new_Sorter100|19181_ ;
  assign \new_Sorter100|19282_  = \new_Sorter100|19182_  & \new_Sorter100|19183_ ;
  assign \new_Sorter100|19283_  = \new_Sorter100|19182_  | \new_Sorter100|19183_ ;
  assign \new_Sorter100|19284_  = \new_Sorter100|19184_  & \new_Sorter100|19185_ ;
  assign \new_Sorter100|19285_  = \new_Sorter100|19184_  | \new_Sorter100|19185_ ;
  assign \new_Sorter100|19286_  = \new_Sorter100|19186_  & \new_Sorter100|19187_ ;
  assign \new_Sorter100|19287_  = \new_Sorter100|19186_  | \new_Sorter100|19187_ ;
  assign \new_Sorter100|19288_  = \new_Sorter100|19188_  & \new_Sorter100|19189_ ;
  assign \new_Sorter100|19289_  = \new_Sorter100|19188_  | \new_Sorter100|19189_ ;
  assign \new_Sorter100|19290_  = \new_Sorter100|19190_  & \new_Sorter100|19191_ ;
  assign \new_Sorter100|19291_  = \new_Sorter100|19190_  | \new_Sorter100|19191_ ;
  assign \new_Sorter100|19292_  = \new_Sorter100|19192_  & \new_Sorter100|19193_ ;
  assign \new_Sorter100|19293_  = \new_Sorter100|19192_  | \new_Sorter100|19193_ ;
  assign \new_Sorter100|19294_  = \new_Sorter100|19194_  & \new_Sorter100|19195_ ;
  assign \new_Sorter100|19295_  = \new_Sorter100|19194_  | \new_Sorter100|19195_ ;
  assign \new_Sorter100|19296_  = \new_Sorter100|19196_  & \new_Sorter100|19197_ ;
  assign \new_Sorter100|19297_  = \new_Sorter100|19196_  | \new_Sorter100|19197_ ;
  assign \new_Sorter100|19298_  = \new_Sorter100|19198_  & \new_Sorter100|19199_ ;
  assign \new_Sorter100|19299_  = \new_Sorter100|19198_  | \new_Sorter100|19199_ ;
  assign \new_Sorter100|19300_  = \new_Sorter100|19200_ ;
  assign \new_Sorter100|19399_  = \new_Sorter100|19299_ ;
  assign \new_Sorter100|19301_  = \new_Sorter100|19201_  & \new_Sorter100|19202_ ;
  assign \new_Sorter100|19302_  = \new_Sorter100|19201_  | \new_Sorter100|19202_ ;
  assign \new_Sorter100|19303_  = \new_Sorter100|19203_  & \new_Sorter100|19204_ ;
  assign \new_Sorter100|19304_  = \new_Sorter100|19203_  | \new_Sorter100|19204_ ;
  assign \new_Sorter100|19305_  = \new_Sorter100|19205_  & \new_Sorter100|19206_ ;
  assign \new_Sorter100|19306_  = \new_Sorter100|19205_  | \new_Sorter100|19206_ ;
  assign \new_Sorter100|19307_  = \new_Sorter100|19207_  & \new_Sorter100|19208_ ;
  assign \new_Sorter100|19308_  = \new_Sorter100|19207_  | \new_Sorter100|19208_ ;
  assign \new_Sorter100|19309_  = \new_Sorter100|19209_  & \new_Sorter100|19210_ ;
  assign \new_Sorter100|19310_  = \new_Sorter100|19209_  | \new_Sorter100|19210_ ;
  assign \new_Sorter100|19311_  = \new_Sorter100|19211_  & \new_Sorter100|19212_ ;
  assign \new_Sorter100|19312_  = \new_Sorter100|19211_  | \new_Sorter100|19212_ ;
  assign \new_Sorter100|19313_  = \new_Sorter100|19213_  & \new_Sorter100|19214_ ;
  assign \new_Sorter100|19314_  = \new_Sorter100|19213_  | \new_Sorter100|19214_ ;
  assign \new_Sorter100|19315_  = \new_Sorter100|19215_  & \new_Sorter100|19216_ ;
  assign \new_Sorter100|19316_  = \new_Sorter100|19215_  | \new_Sorter100|19216_ ;
  assign \new_Sorter100|19317_  = \new_Sorter100|19217_  & \new_Sorter100|19218_ ;
  assign \new_Sorter100|19318_  = \new_Sorter100|19217_  | \new_Sorter100|19218_ ;
  assign \new_Sorter100|19319_  = \new_Sorter100|19219_  & \new_Sorter100|19220_ ;
  assign \new_Sorter100|19320_  = \new_Sorter100|19219_  | \new_Sorter100|19220_ ;
  assign \new_Sorter100|19321_  = \new_Sorter100|19221_  & \new_Sorter100|19222_ ;
  assign \new_Sorter100|19322_  = \new_Sorter100|19221_  | \new_Sorter100|19222_ ;
  assign \new_Sorter100|19323_  = \new_Sorter100|19223_  & \new_Sorter100|19224_ ;
  assign \new_Sorter100|19324_  = \new_Sorter100|19223_  | \new_Sorter100|19224_ ;
  assign \new_Sorter100|19325_  = \new_Sorter100|19225_  & \new_Sorter100|19226_ ;
  assign \new_Sorter100|19326_  = \new_Sorter100|19225_  | \new_Sorter100|19226_ ;
  assign \new_Sorter100|19327_  = \new_Sorter100|19227_  & \new_Sorter100|19228_ ;
  assign \new_Sorter100|19328_  = \new_Sorter100|19227_  | \new_Sorter100|19228_ ;
  assign \new_Sorter100|19329_  = \new_Sorter100|19229_  & \new_Sorter100|19230_ ;
  assign \new_Sorter100|19330_  = \new_Sorter100|19229_  | \new_Sorter100|19230_ ;
  assign \new_Sorter100|19331_  = \new_Sorter100|19231_  & \new_Sorter100|19232_ ;
  assign \new_Sorter100|19332_  = \new_Sorter100|19231_  | \new_Sorter100|19232_ ;
  assign \new_Sorter100|19333_  = \new_Sorter100|19233_  & \new_Sorter100|19234_ ;
  assign \new_Sorter100|19334_  = \new_Sorter100|19233_  | \new_Sorter100|19234_ ;
  assign \new_Sorter100|19335_  = \new_Sorter100|19235_  & \new_Sorter100|19236_ ;
  assign \new_Sorter100|19336_  = \new_Sorter100|19235_  | \new_Sorter100|19236_ ;
  assign \new_Sorter100|19337_  = \new_Sorter100|19237_  & \new_Sorter100|19238_ ;
  assign \new_Sorter100|19338_  = \new_Sorter100|19237_  | \new_Sorter100|19238_ ;
  assign \new_Sorter100|19339_  = \new_Sorter100|19239_  & \new_Sorter100|19240_ ;
  assign \new_Sorter100|19340_  = \new_Sorter100|19239_  | \new_Sorter100|19240_ ;
  assign \new_Sorter100|19341_  = \new_Sorter100|19241_  & \new_Sorter100|19242_ ;
  assign \new_Sorter100|19342_  = \new_Sorter100|19241_  | \new_Sorter100|19242_ ;
  assign \new_Sorter100|19343_  = \new_Sorter100|19243_  & \new_Sorter100|19244_ ;
  assign \new_Sorter100|19344_  = \new_Sorter100|19243_  | \new_Sorter100|19244_ ;
  assign \new_Sorter100|19345_  = \new_Sorter100|19245_  & \new_Sorter100|19246_ ;
  assign \new_Sorter100|19346_  = \new_Sorter100|19245_  | \new_Sorter100|19246_ ;
  assign \new_Sorter100|19347_  = \new_Sorter100|19247_  & \new_Sorter100|19248_ ;
  assign \new_Sorter100|19348_  = \new_Sorter100|19247_  | \new_Sorter100|19248_ ;
  assign \new_Sorter100|19349_  = \new_Sorter100|19249_  & \new_Sorter100|19250_ ;
  assign \new_Sorter100|19350_  = \new_Sorter100|19249_  | \new_Sorter100|19250_ ;
  assign \new_Sorter100|19351_  = \new_Sorter100|19251_  & \new_Sorter100|19252_ ;
  assign \new_Sorter100|19352_  = \new_Sorter100|19251_  | \new_Sorter100|19252_ ;
  assign \new_Sorter100|19353_  = \new_Sorter100|19253_  & \new_Sorter100|19254_ ;
  assign \new_Sorter100|19354_  = \new_Sorter100|19253_  | \new_Sorter100|19254_ ;
  assign \new_Sorter100|19355_  = \new_Sorter100|19255_  & \new_Sorter100|19256_ ;
  assign \new_Sorter100|19356_  = \new_Sorter100|19255_  | \new_Sorter100|19256_ ;
  assign \new_Sorter100|19357_  = \new_Sorter100|19257_  & \new_Sorter100|19258_ ;
  assign \new_Sorter100|19358_  = \new_Sorter100|19257_  | \new_Sorter100|19258_ ;
  assign \new_Sorter100|19359_  = \new_Sorter100|19259_  & \new_Sorter100|19260_ ;
  assign \new_Sorter100|19360_  = \new_Sorter100|19259_  | \new_Sorter100|19260_ ;
  assign \new_Sorter100|19361_  = \new_Sorter100|19261_  & \new_Sorter100|19262_ ;
  assign \new_Sorter100|19362_  = \new_Sorter100|19261_  | \new_Sorter100|19262_ ;
  assign \new_Sorter100|19363_  = \new_Sorter100|19263_  & \new_Sorter100|19264_ ;
  assign \new_Sorter100|19364_  = \new_Sorter100|19263_  | \new_Sorter100|19264_ ;
  assign \new_Sorter100|19365_  = \new_Sorter100|19265_  & \new_Sorter100|19266_ ;
  assign \new_Sorter100|19366_  = \new_Sorter100|19265_  | \new_Sorter100|19266_ ;
  assign \new_Sorter100|19367_  = \new_Sorter100|19267_  & \new_Sorter100|19268_ ;
  assign \new_Sorter100|19368_  = \new_Sorter100|19267_  | \new_Sorter100|19268_ ;
  assign \new_Sorter100|19369_  = \new_Sorter100|19269_  & \new_Sorter100|19270_ ;
  assign \new_Sorter100|19370_  = \new_Sorter100|19269_  | \new_Sorter100|19270_ ;
  assign \new_Sorter100|19371_  = \new_Sorter100|19271_  & \new_Sorter100|19272_ ;
  assign \new_Sorter100|19372_  = \new_Sorter100|19271_  | \new_Sorter100|19272_ ;
  assign \new_Sorter100|19373_  = \new_Sorter100|19273_  & \new_Sorter100|19274_ ;
  assign \new_Sorter100|19374_  = \new_Sorter100|19273_  | \new_Sorter100|19274_ ;
  assign \new_Sorter100|19375_  = \new_Sorter100|19275_  & \new_Sorter100|19276_ ;
  assign \new_Sorter100|19376_  = \new_Sorter100|19275_  | \new_Sorter100|19276_ ;
  assign \new_Sorter100|19377_  = \new_Sorter100|19277_  & \new_Sorter100|19278_ ;
  assign \new_Sorter100|19378_  = \new_Sorter100|19277_  | \new_Sorter100|19278_ ;
  assign \new_Sorter100|19379_  = \new_Sorter100|19279_  & \new_Sorter100|19280_ ;
  assign \new_Sorter100|19380_  = \new_Sorter100|19279_  | \new_Sorter100|19280_ ;
  assign \new_Sorter100|19381_  = \new_Sorter100|19281_  & \new_Sorter100|19282_ ;
  assign \new_Sorter100|19382_  = \new_Sorter100|19281_  | \new_Sorter100|19282_ ;
  assign \new_Sorter100|19383_  = \new_Sorter100|19283_  & \new_Sorter100|19284_ ;
  assign \new_Sorter100|19384_  = \new_Sorter100|19283_  | \new_Sorter100|19284_ ;
  assign \new_Sorter100|19385_  = \new_Sorter100|19285_  & \new_Sorter100|19286_ ;
  assign \new_Sorter100|19386_  = \new_Sorter100|19285_  | \new_Sorter100|19286_ ;
  assign \new_Sorter100|19387_  = \new_Sorter100|19287_  & \new_Sorter100|19288_ ;
  assign \new_Sorter100|19388_  = \new_Sorter100|19287_  | \new_Sorter100|19288_ ;
  assign \new_Sorter100|19389_  = \new_Sorter100|19289_  & \new_Sorter100|19290_ ;
  assign \new_Sorter100|19390_  = \new_Sorter100|19289_  | \new_Sorter100|19290_ ;
  assign \new_Sorter100|19391_  = \new_Sorter100|19291_  & \new_Sorter100|19292_ ;
  assign \new_Sorter100|19392_  = \new_Sorter100|19291_  | \new_Sorter100|19292_ ;
  assign \new_Sorter100|19393_  = \new_Sorter100|19293_  & \new_Sorter100|19294_ ;
  assign \new_Sorter100|19394_  = \new_Sorter100|19293_  | \new_Sorter100|19294_ ;
  assign \new_Sorter100|19395_  = \new_Sorter100|19295_  & \new_Sorter100|19296_ ;
  assign \new_Sorter100|19396_  = \new_Sorter100|19295_  | \new_Sorter100|19296_ ;
  assign \new_Sorter100|19397_  = \new_Sorter100|19297_  & \new_Sorter100|19298_ ;
  assign \new_Sorter100|19398_  = \new_Sorter100|19297_  | \new_Sorter100|19298_ ;
  assign \new_Sorter100|19400_  = \new_Sorter100|19300_  & \new_Sorter100|19301_ ;
  assign \new_Sorter100|19401_  = \new_Sorter100|19300_  | \new_Sorter100|19301_ ;
  assign \new_Sorter100|19402_  = \new_Sorter100|19302_  & \new_Sorter100|19303_ ;
  assign \new_Sorter100|19403_  = \new_Sorter100|19302_  | \new_Sorter100|19303_ ;
  assign \new_Sorter100|19404_  = \new_Sorter100|19304_  & \new_Sorter100|19305_ ;
  assign \new_Sorter100|19405_  = \new_Sorter100|19304_  | \new_Sorter100|19305_ ;
  assign \new_Sorter100|19406_  = \new_Sorter100|19306_  & \new_Sorter100|19307_ ;
  assign \new_Sorter100|19407_  = \new_Sorter100|19306_  | \new_Sorter100|19307_ ;
  assign \new_Sorter100|19408_  = \new_Sorter100|19308_  & \new_Sorter100|19309_ ;
  assign \new_Sorter100|19409_  = \new_Sorter100|19308_  | \new_Sorter100|19309_ ;
  assign \new_Sorter100|19410_  = \new_Sorter100|19310_  & \new_Sorter100|19311_ ;
  assign \new_Sorter100|19411_  = \new_Sorter100|19310_  | \new_Sorter100|19311_ ;
  assign \new_Sorter100|19412_  = \new_Sorter100|19312_  & \new_Sorter100|19313_ ;
  assign \new_Sorter100|19413_  = \new_Sorter100|19312_  | \new_Sorter100|19313_ ;
  assign \new_Sorter100|19414_  = \new_Sorter100|19314_  & \new_Sorter100|19315_ ;
  assign \new_Sorter100|19415_  = \new_Sorter100|19314_  | \new_Sorter100|19315_ ;
  assign \new_Sorter100|19416_  = \new_Sorter100|19316_  & \new_Sorter100|19317_ ;
  assign \new_Sorter100|19417_  = \new_Sorter100|19316_  | \new_Sorter100|19317_ ;
  assign \new_Sorter100|19418_  = \new_Sorter100|19318_  & \new_Sorter100|19319_ ;
  assign \new_Sorter100|19419_  = \new_Sorter100|19318_  | \new_Sorter100|19319_ ;
  assign \new_Sorter100|19420_  = \new_Sorter100|19320_  & \new_Sorter100|19321_ ;
  assign \new_Sorter100|19421_  = \new_Sorter100|19320_  | \new_Sorter100|19321_ ;
  assign \new_Sorter100|19422_  = \new_Sorter100|19322_  & \new_Sorter100|19323_ ;
  assign \new_Sorter100|19423_  = \new_Sorter100|19322_  | \new_Sorter100|19323_ ;
  assign \new_Sorter100|19424_  = \new_Sorter100|19324_  & \new_Sorter100|19325_ ;
  assign \new_Sorter100|19425_  = \new_Sorter100|19324_  | \new_Sorter100|19325_ ;
  assign \new_Sorter100|19426_  = \new_Sorter100|19326_  & \new_Sorter100|19327_ ;
  assign \new_Sorter100|19427_  = \new_Sorter100|19326_  | \new_Sorter100|19327_ ;
  assign \new_Sorter100|19428_  = \new_Sorter100|19328_  & \new_Sorter100|19329_ ;
  assign \new_Sorter100|19429_  = \new_Sorter100|19328_  | \new_Sorter100|19329_ ;
  assign \new_Sorter100|19430_  = \new_Sorter100|19330_  & \new_Sorter100|19331_ ;
  assign \new_Sorter100|19431_  = \new_Sorter100|19330_  | \new_Sorter100|19331_ ;
  assign \new_Sorter100|19432_  = \new_Sorter100|19332_  & \new_Sorter100|19333_ ;
  assign \new_Sorter100|19433_  = \new_Sorter100|19332_  | \new_Sorter100|19333_ ;
  assign \new_Sorter100|19434_  = \new_Sorter100|19334_  & \new_Sorter100|19335_ ;
  assign \new_Sorter100|19435_  = \new_Sorter100|19334_  | \new_Sorter100|19335_ ;
  assign \new_Sorter100|19436_  = \new_Sorter100|19336_  & \new_Sorter100|19337_ ;
  assign \new_Sorter100|19437_  = \new_Sorter100|19336_  | \new_Sorter100|19337_ ;
  assign \new_Sorter100|19438_  = \new_Sorter100|19338_  & \new_Sorter100|19339_ ;
  assign \new_Sorter100|19439_  = \new_Sorter100|19338_  | \new_Sorter100|19339_ ;
  assign \new_Sorter100|19440_  = \new_Sorter100|19340_  & \new_Sorter100|19341_ ;
  assign \new_Sorter100|19441_  = \new_Sorter100|19340_  | \new_Sorter100|19341_ ;
  assign \new_Sorter100|19442_  = \new_Sorter100|19342_  & \new_Sorter100|19343_ ;
  assign \new_Sorter100|19443_  = \new_Sorter100|19342_  | \new_Sorter100|19343_ ;
  assign \new_Sorter100|19444_  = \new_Sorter100|19344_  & \new_Sorter100|19345_ ;
  assign \new_Sorter100|19445_  = \new_Sorter100|19344_  | \new_Sorter100|19345_ ;
  assign \new_Sorter100|19446_  = \new_Sorter100|19346_  & \new_Sorter100|19347_ ;
  assign \new_Sorter100|19447_  = \new_Sorter100|19346_  | \new_Sorter100|19347_ ;
  assign \new_Sorter100|19448_  = \new_Sorter100|19348_  & \new_Sorter100|19349_ ;
  assign \new_Sorter100|19449_  = \new_Sorter100|19348_  | \new_Sorter100|19349_ ;
  assign \new_Sorter100|19450_  = \new_Sorter100|19350_  & \new_Sorter100|19351_ ;
  assign \new_Sorter100|19451_  = \new_Sorter100|19350_  | \new_Sorter100|19351_ ;
  assign \new_Sorter100|19452_  = \new_Sorter100|19352_  & \new_Sorter100|19353_ ;
  assign \new_Sorter100|19453_  = \new_Sorter100|19352_  | \new_Sorter100|19353_ ;
  assign \new_Sorter100|19454_  = \new_Sorter100|19354_  & \new_Sorter100|19355_ ;
  assign \new_Sorter100|19455_  = \new_Sorter100|19354_  | \new_Sorter100|19355_ ;
  assign \new_Sorter100|19456_  = \new_Sorter100|19356_  & \new_Sorter100|19357_ ;
  assign \new_Sorter100|19457_  = \new_Sorter100|19356_  | \new_Sorter100|19357_ ;
  assign \new_Sorter100|19458_  = \new_Sorter100|19358_  & \new_Sorter100|19359_ ;
  assign \new_Sorter100|19459_  = \new_Sorter100|19358_  | \new_Sorter100|19359_ ;
  assign \new_Sorter100|19460_  = \new_Sorter100|19360_  & \new_Sorter100|19361_ ;
  assign \new_Sorter100|19461_  = \new_Sorter100|19360_  | \new_Sorter100|19361_ ;
  assign \new_Sorter100|19462_  = \new_Sorter100|19362_  & \new_Sorter100|19363_ ;
  assign \new_Sorter100|19463_  = \new_Sorter100|19362_  | \new_Sorter100|19363_ ;
  assign \new_Sorter100|19464_  = \new_Sorter100|19364_  & \new_Sorter100|19365_ ;
  assign \new_Sorter100|19465_  = \new_Sorter100|19364_  | \new_Sorter100|19365_ ;
  assign \new_Sorter100|19466_  = \new_Sorter100|19366_  & \new_Sorter100|19367_ ;
  assign \new_Sorter100|19467_  = \new_Sorter100|19366_  | \new_Sorter100|19367_ ;
  assign \new_Sorter100|19468_  = \new_Sorter100|19368_  & \new_Sorter100|19369_ ;
  assign \new_Sorter100|19469_  = \new_Sorter100|19368_  | \new_Sorter100|19369_ ;
  assign \new_Sorter100|19470_  = \new_Sorter100|19370_  & \new_Sorter100|19371_ ;
  assign \new_Sorter100|19471_  = \new_Sorter100|19370_  | \new_Sorter100|19371_ ;
  assign \new_Sorter100|19472_  = \new_Sorter100|19372_  & \new_Sorter100|19373_ ;
  assign \new_Sorter100|19473_  = \new_Sorter100|19372_  | \new_Sorter100|19373_ ;
  assign \new_Sorter100|19474_  = \new_Sorter100|19374_  & \new_Sorter100|19375_ ;
  assign \new_Sorter100|19475_  = \new_Sorter100|19374_  | \new_Sorter100|19375_ ;
  assign \new_Sorter100|19476_  = \new_Sorter100|19376_  & \new_Sorter100|19377_ ;
  assign \new_Sorter100|19477_  = \new_Sorter100|19376_  | \new_Sorter100|19377_ ;
  assign \new_Sorter100|19478_  = \new_Sorter100|19378_  & \new_Sorter100|19379_ ;
  assign \new_Sorter100|19479_  = \new_Sorter100|19378_  | \new_Sorter100|19379_ ;
  assign \new_Sorter100|19480_  = \new_Sorter100|19380_  & \new_Sorter100|19381_ ;
  assign \new_Sorter100|19481_  = \new_Sorter100|19380_  | \new_Sorter100|19381_ ;
  assign \new_Sorter100|19482_  = \new_Sorter100|19382_  & \new_Sorter100|19383_ ;
  assign \new_Sorter100|19483_  = \new_Sorter100|19382_  | \new_Sorter100|19383_ ;
  assign \new_Sorter100|19484_  = \new_Sorter100|19384_  & \new_Sorter100|19385_ ;
  assign \new_Sorter100|19485_  = \new_Sorter100|19384_  | \new_Sorter100|19385_ ;
  assign \new_Sorter100|19486_  = \new_Sorter100|19386_  & \new_Sorter100|19387_ ;
  assign \new_Sorter100|19487_  = \new_Sorter100|19386_  | \new_Sorter100|19387_ ;
  assign \new_Sorter100|19488_  = \new_Sorter100|19388_  & \new_Sorter100|19389_ ;
  assign \new_Sorter100|19489_  = \new_Sorter100|19388_  | \new_Sorter100|19389_ ;
  assign \new_Sorter100|19490_  = \new_Sorter100|19390_  & \new_Sorter100|19391_ ;
  assign \new_Sorter100|19491_  = \new_Sorter100|19390_  | \new_Sorter100|19391_ ;
  assign \new_Sorter100|19492_  = \new_Sorter100|19392_  & \new_Sorter100|19393_ ;
  assign \new_Sorter100|19493_  = \new_Sorter100|19392_  | \new_Sorter100|19393_ ;
  assign \new_Sorter100|19494_  = \new_Sorter100|19394_  & \new_Sorter100|19395_ ;
  assign \new_Sorter100|19495_  = \new_Sorter100|19394_  | \new_Sorter100|19395_ ;
  assign \new_Sorter100|19496_  = \new_Sorter100|19396_  & \new_Sorter100|19397_ ;
  assign \new_Sorter100|19497_  = \new_Sorter100|19396_  | \new_Sorter100|19397_ ;
  assign \new_Sorter100|19498_  = \new_Sorter100|19398_  & \new_Sorter100|19399_ ;
  assign \new_Sorter100|19499_  = \new_Sorter100|19398_  | \new_Sorter100|19399_ ;
  assign \new_Sorter100|19500_  = \new_Sorter100|19400_ ;
  assign \new_Sorter100|19599_  = \new_Sorter100|19499_ ;
  assign \new_Sorter100|19501_  = \new_Sorter100|19401_  & \new_Sorter100|19402_ ;
  assign \new_Sorter100|19502_  = \new_Sorter100|19401_  | \new_Sorter100|19402_ ;
  assign \new_Sorter100|19503_  = \new_Sorter100|19403_  & \new_Sorter100|19404_ ;
  assign \new_Sorter100|19504_  = \new_Sorter100|19403_  | \new_Sorter100|19404_ ;
  assign \new_Sorter100|19505_  = \new_Sorter100|19405_  & \new_Sorter100|19406_ ;
  assign \new_Sorter100|19506_  = \new_Sorter100|19405_  | \new_Sorter100|19406_ ;
  assign \new_Sorter100|19507_  = \new_Sorter100|19407_  & \new_Sorter100|19408_ ;
  assign \new_Sorter100|19508_  = \new_Sorter100|19407_  | \new_Sorter100|19408_ ;
  assign \new_Sorter100|19509_  = \new_Sorter100|19409_  & \new_Sorter100|19410_ ;
  assign \new_Sorter100|19510_  = \new_Sorter100|19409_  | \new_Sorter100|19410_ ;
  assign \new_Sorter100|19511_  = \new_Sorter100|19411_  & \new_Sorter100|19412_ ;
  assign \new_Sorter100|19512_  = \new_Sorter100|19411_  | \new_Sorter100|19412_ ;
  assign \new_Sorter100|19513_  = \new_Sorter100|19413_  & \new_Sorter100|19414_ ;
  assign \new_Sorter100|19514_  = \new_Sorter100|19413_  | \new_Sorter100|19414_ ;
  assign \new_Sorter100|19515_  = \new_Sorter100|19415_  & \new_Sorter100|19416_ ;
  assign \new_Sorter100|19516_  = \new_Sorter100|19415_  | \new_Sorter100|19416_ ;
  assign \new_Sorter100|19517_  = \new_Sorter100|19417_  & \new_Sorter100|19418_ ;
  assign \new_Sorter100|19518_  = \new_Sorter100|19417_  | \new_Sorter100|19418_ ;
  assign \new_Sorter100|19519_  = \new_Sorter100|19419_  & \new_Sorter100|19420_ ;
  assign \new_Sorter100|19520_  = \new_Sorter100|19419_  | \new_Sorter100|19420_ ;
  assign \new_Sorter100|19521_  = \new_Sorter100|19421_  & \new_Sorter100|19422_ ;
  assign \new_Sorter100|19522_  = \new_Sorter100|19421_  | \new_Sorter100|19422_ ;
  assign \new_Sorter100|19523_  = \new_Sorter100|19423_  & \new_Sorter100|19424_ ;
  assign \new_Sorter100|19524_  = \new_Sorter100|19423_  | \new_Sorter100|19424_ ;
  assign \new_Sorter100|19525_  = \new_Sorter100|19425_  & \new_Sorter100|19426_ ;
  assign \new_Sorter100|19526_  = \new_Sorter100|19425_  | \new_Sorter100|19426_ ;
  assign \new_Sorter100|19527_  = \new_Sorter100|19427_  & \new_Sorter100|19428_ ;
  assign \new_Sorter100|19528_  = \new_Sorter100|19427_  | \new_Sorter100|19428_ ;
  assign \new_Sorter100|19529_  = \new_Sorter100|19429_  & \new_Sorter100|19430_ ;
  assign \new_Sorter100|19530_  = \new_Sorter100|19429_  | \new_Sorter100|19430_ ;
  assign \new_Sorter100|19531_  = \new_Sorter100|19431_  & \new_Sorter100|19432_ ;
  assign \new_Sorter100|19532_  = \new_Sorter100|19431_  | \new_Sorter100|19432_ ;
  assign \new_Sorter100|19533_  = \new_Sorter100|19433_  & \new_Sorter100|19434_ ;
  assign \new_Sorter100|19534_  = \new_Sorter100|19433_  | \new_Sorter100|19434_ ;
  assign \new_Sorter100|19535_  = \new_Sorter100|19435_  & \new_Sorter100|19436_ ;
  assign \new_Sorter100|19536_  = \new_Sorter100|19435_  | \new_Sorter100|19436_ ;
  assign \new_Sorter100|19537_  = \new_Sorter100|19437_  & \new_Sorter100|19438_ ;
  assign \new_Sorter100|19538_  = \new_Sorter100|19437_  | \new_Sorter100|19438_ ;
  assign \new_Sorter100|19539_  = \new_Sorter100|19439_  & \new_Sorter100|19440_ ;
  assign \new_Sorter100|19540_  = \new_Sorter100|19439_  | \new_Sorter100|19440_ ;
  assign \new_Sorter100|19541_  = \new_Sorter100|19441_  & \new_Sorter100|19442_ ;
  assign \new_Sorter100|19542_  = \new_Sorter100|19441_  | \new_Sorter100|19442_ ;
  assign \new_Sorter100|19543_  = \new_Sorter100|19443_  & \new_Sorter100|19444_ ;
  assign \new_Sorter100|19544_  = \new_Sorter100|19443_  | \new_Sorter100|19444_ ;
  assign \new_Sorter100|19545_  = \new_Sorter100|19445_  & \new_Sorter100|19446_ ;
  assign \new_Sorter100|19546_  = \new_Sorter100|19445_  | \new_Sorter100|19446_ ;
  assign \new_Sorter100|19547_  = \new_Sorter100|19447_  & \new_Sorter100|19448_ ;
  assign \new_Sorter100|19548_  = \new_Sorter100|19447_  | \new_Sorter100|19448_ ;
  assign \new_Sorter100|19549_  = \new_Sorter100|19449_  & \new_Sorter100|19450_ ;
  assign \new_Sorter100|19550_  = \new_Sorter100|19449_  | \new_Sorter100|19450_ ;
  assign \new_Sorter100|19551_  = \new_Sorter100|19451_  & \new_Sorter100|19452_ ;
  assign \new_Sorter100|19552_  = \new_Sorter100|19451_  | \new_Sorter100|19452_ ;
  assign \new_Sorter100|19553_  = \new_Sorter100|19453_  & \new_Sorter100|19454_ ;
  assign \new_Sorter100|19554_  = \new_Sorter100|19453_  | \new_Sorter100|19454_ ;
  assign \new_Sorter100|19555_  = \new_Sorter100|19455_  & \new_Sorter100|19456_ ;
  assign \new_Sorter100|19556_  = \new_Sorter100|19455_  | \new_Sorter100|19456_ ;
  assign \new_Sorter100|19557_  = \new_Sorter100|19457_  & \new_Sorter100|19458_ ;
  assign \new_Sorter100|19558_  = \new_Sorter100|19457_  | \new_Sorter100|19458_ ;
  assign \new_Sorter100|19559_  = \new_Sorter100|19459_  & \new_Sorter100|19460_ ;
  assign \new_Sorter100|19560_  = \new_Sorter100|19459_  | \new_Sorter100|19460_ ;
  assign \new_Sorter100|19561_  = \new_Sorter100|19461_  & \new_Sorter100|19462_ ;
  assign \new_Sorter100|19562_  = \new_Sorter100|19461_  | \new_Sorter100|19462_ ;
  assign \new_Sorter100|19563_  = \new_Sorter100|19463_  & \new_Sorter100|19464_ ;
  assign \new_Sorter100|19564_  = \new_Sorter100|19463_  | \new_Sorter100|19464_ ;
  assign \new_Sorter100|19565_  = \new_Sorter100|19465_  & \new_Sorter100|19466_ ;
  assign \new_Sorter100|19566_  = \new_Sorter100|19465_  | \new_Sorter100|19466_ ;
  assign \new_Sorter100|19567_  = \new_Sorter100|19467_  & \new_Sorter100|19468_ ;
  assign \new_Sorter100|19568_  = \new_Sorter100|19467_  | \new_Sorter100|19468_ ;
  assign \new_Sorter100|19569_  = \new_Sorter100|19469_  & \new_Sorter100|19470_ ;
  assign \new_Sorter100|19570_  = \new_Sorter100|19469_  | \new_Sorter100|19470_ ;
  assign \new_Sorter100|19571_  = \new_Sorter100|19471_  & \new_Sorter100|19472_ ;
  assign \new_Sorter100|19572_  = \new_Sorter100|19471_  | \new_Sorter100|19472_ ;
  assign \new_Sorter100|19573_  = \new_Sorter100|19473_  & \new_Sorter100|19474_ ;
  assign \new_Sorter100|19574_  = \new_Sorter100|19473_  | \new_Sorter100|19474_ ;
  assign \new_Sorter100|19575_  = \new_Sorter100|19475_  & \new_Sorter100|19476_ ;
  assign \new_Sorter100|19576_  = \new_Sorter100|19475_  | \new_Sorter100|19476_ ;
  assign \new_Sorter100|19577_  = \new_Sorter100|19477_  & \new_Sorter100|19478_ ;
  assign \new_Sorter100|19578_  = \new_Sorter100|19477_  | \new_Sorter100|19478_ ;
  assign \new_Sorter100|19579_  = \new_Sorter100|19479_  & \new_Sorter100|19480_ ;
  assign \new_Sorter100|19580_  = \new_Sorter100|19479_  | \new_Sorter100|19480_ ;
  assign \new_Sorter100|19581_  = \new_Sorter100|19481_  & \new_Sorter100|19482_ ;
  assign \new_Sorter100|19582_  = \new_Sorter100|19481_  | \new_Sorter100|19482_ ;
  assign \new_Sorter100|19583_  = \new_Sorter100|19483_  & \new_Sorter100|19484_ ;
  assign \new_Sorter100|19584_  = \new_Sorter100|19483_  | \new_Sorter100|19484_ ;
  assign \new_Sorter100|19585_  = \new_Sorter100|19485_  & \new_Sorter100|19486_ ;
  assign \new_Sorter100|19586_  = \new_Sorter100|19485_  | \new_Sorter100|19486_ ;
  assign \new_Sorter100|19587_  = \new_Sorter100|19487_  & \new_Sorter100|19488_ ;
  assign \new_Sorter100|19588_  = \new_Sorter100|19487_  | \new_Sorter100|19488_ ;
  assign \new_Sorter100|19589_  = \new_Sorter100|19489_  & \new_Sorter100|19490_ ;
  assign \new_Sorter100|19590_  = \new_Sorter100|19489_  | \new_Sorter100|19490_ ;
  assign \new_Sorter100|19591_  = \new_Sorter100|19491_  & \new_Sorter100|19492_ ;
  assign \new_Sorter100|19592_  = \new_Sorter100|19491_  | \new_Sorter100|19492_ ;
  assign \new_Sorter100|19593_  = \new_Sorter100|19493_  & \new_Sorter100|19494_ ;
  assign \new_Sorter100|19594_  = \new_Sorter100|19493_  | \new_Sorter100|19494_ ;
  assign \new_Sorter100|19595_  = \new_Sorter100|19495_  & \new_Sorter100|19496_ ;
  assign \new_Sorter100|19596_  = \new_Sorter100|19495_  | \new_Sorter100|19496_ ;
  assign \new_Sorter100|19597_  = \new_Sorter100|19497_  & \new_Sorter100|19498_ ;
  assign \new_Sorter100|19598_  = \new_Sorter100|19497_  | \new_Sorter100|19498_ ;
  assign \new_Sorter100|19600_  = \new_Sorter100|19500_  & \new_Sorter100|19501_ ;
  assign \new_Sorter100|19601_  = \new_Sorter100|19500_  | \new_Sorter100|19501_ ;
  assign \new_Sorter100|19602_  = \new_Sorter100|19502_  & \new_Sorter100|19503_ ;
  assign \new_Sorter100|19603_  = \new_Sorter100|19502_  | \new_Sorter100|19503_ ;
  assign \new_Sorter100|19604_  = \new_Sorter100|19504_  & \new_Sorter100|19505_ ;
  assign \new_Sorter100|19605_  = \new_Sorter100|19504_  | \new_Sorter100|19505_ ;
  assign \new_Sorter100|19606_  = \new_Sorter100|19506_  & \new_Sorter100|19507_ ;
  assign \new_Sorter100|19607_  = \new_Sorter100|19506_  | \new_Sorter100|19507_ ;
  assign \new_Sorter100|19608_  = \new_Sorter100|19508_  & \new_Sorter100|19509_ ;
  assign \new_Sorter100|19609_  = \new_Sorter100|19508_  | \new_Sorter100|19509_ ;
  assign \new_Sorter100|19610_  = \new_Sorter100|19510_  & \new_Sorter100|19511_ ;
  assign \new_Sorter100|19611_  = \new_Sorter100|19510_  | \new_Sorter100|19511_ ;
  assign \new_Sorter100|19612_  = \new_Sorter100|19512_  & \new_Sorter100|19513_ ;
  assign \new_Sorter100|19613_  = \new_Sorter100|19512_  | \new_Sorter100|19513_ ;
  assign \new_Sorter100|19614_  = \new_Sorter100|19514_  & \new_Sorter100|19515_ ;
  assign \new_Sorter100|19615_  = \new_Sorter100|19514_  | \new_Sorter100|19515_ ;
  assign \new_Sorter100|19616_  = \new_Sorter100|19516_  & \new_Sorter100|19517_ ;
  assign \new_Sorter100|19617_  = \new_Sorter100|19516_  | \new_Sorter100|19517_ ;
  assign \new_Sorter100|19618_  = \new_Sorter100|19518_  & \new_Sorter100|19519_ ;
  assign \new_Sorter100|19619_  = \new_Sorter100|19518_  | \new_Sorter100|19519_ ;
  assign \new_Sorter100|19620_  = \new_Sorter100|19520_  & \new_Sorter100|19521_ ;
  assign \new_Sorter100|19621_  = \new_Sorter100|19520_  | \new_Sorter100|19521_ ;
  assign \new_Sorter100|19622_  = \new_Sorter100|19522_  & \new_Sorter100|19523_ ;
  assign \new_Sorter100|19623_  = \new_Sorter100|19522_  | \new_Sorter100|19523_ ;
  assign \new_Sorter100|19624_  = \new_Sorter100|19524_  & \new_Sorter100|19525_ ;
  assign \new_Sorter100|19625_  = \new_Sorter100|19524_  | \new_Sorter100|19525_ ;
  assign \new_Sorter100|19626_  = \new_Sorter100|19526_  & \new_Sorter100|19527_ ;
  assign \new_Sorter100|19627_  = \new_Sorter100|19526_  | \new_Sorter100|19527_ ;
  assign \new_Sorter100|19628_  = \new_Sorter100|19528_  & \new_Sorter100|19529_ ;
  assign \new_Sorter100|19629_  = \new_Sorter100|19528_  | \new_Sorter100|19529_ ;
  assign \new_Sorter100|19630_  = \new_Sorter100|19530_  & \new_Sorter100|19531_ ;
  assign \new_Sorter100|19631_  = \new_Sorter100|19530_  | \new_Sorter100|19531_ ;
  assign \new_Sorter100|19632_  = \new_Sorter100|19532_  & \new_Sorter100|19533_ ;
  assign \new_Sorter100|19633_  = \new_Sorter100|19532_  | \new_Sorter100|19533_ ;
  assign \new_Sorter100|19634_  = \new_Sorter100|19534_  & \new_Sorter100|19535_ ;
  assign \new_Sorter100|19635_  = \new_Sorter100|19534_  | \new_Sorter100|19535_ ;
  assign \new_Sorter100|19636_  = \new_Sorter100|19536_  & \new_Sorter100|19537_ ;
  assign \new_Sorter100|19637_  = \new_Sorter100|19536_  | \new_Sorter100|19537_ ;
  assign \new_Sorter100|19638_  = \new_Sorter100|19538_  & \new_Sorter100|19539_ ;
  assign \new_Sorter100|19639_  = \new_Sorter100|19538_  | \new_Sorter100|19539_ ;
  assign \new_Sorter100|19640_  = \new_Sorter100|19540_  & \new_Sorter100|19541_ ;
  assign \new_Sorter100|19641_  = \new_Sorter100|19540_  | \new_Sorter100|19541_ ;
  assign \new_Sorter100|19642_  = \new_Sorter100|19542_  & \new_Sorter100|19543_ ;
  assign \new_Sorter100|19643_  = \new_Sorter100|19542_  | \new_Sorter100|19543_ ;
  assign \new_Sorter100|19644_  = \new_Sorter100|19544_  & \new_Sorter100|19545_ ;
  assign \new_Sorter100|19645_  = \new_Sorter100|19544_  | \new_Sorter100|19545_ ;
  assign \new_Sorter100|19646_  = \new_Sorter100|19546_  & \new_Sorter100|19547_ ;
  assign \new_Sorter100|19647_  = \new_Sorter100|19546_  | \new_Sorter100|19547_ ;
  assign \new_Sorter100|19648_  = \new_Sorter100|19548_  & \new_Sorter100|19549_ ;
  assign \new_Sorter100|19649_  = \new_Sorter100|19548_  | \new_Sorter100|19549_ ;
  assign \new_Sorter100|19650_  = \new_Sorter100|19550_  & \new_Sorter100|19551_ ;
  assign \new_Sorter100|19651_  = \new_Sorter100|19550_  | \new_Sorter100|19551_ ;
  assign \new_Sorter100|19652_  = \new_Sorter100|19552_  & \new_Sorter100|19553_ ;
  assign \new_Sorter100|19653_  = \new_Sorter100|19552_  | \new_Sorter100|19553_ ;
  assign \new_Sorter100|19654_  = \new_Sorter100|19554_  & \new_Sorter100|19555_ ;
  assign \new_Sorter100|19655_  = \new_Sorter100|19554_  | \new_Sorter100|19555_ ;
  assign \new_Sorter100|19656_  = \new_Sorter100|19556_  & \new_Sorter100|19557_ ;
  assign \new_Sorter100|19657_  = \new_Sorter100|19556_  | \new_Sorter100|19557_ ;
  assign \new_Sorter100|19658_  = \new_Sorter100|19558_  & \new_Sorter100|19559_ ;
  assign \new_Sorter100|19659_  = \new_Sorter100|19558_  | \new_Sorter100|19559_ ;
  assign \new_Sorter100|19660_  = \new_Sorter100|19560_  & \new_Sorter100|19561_ ;
  assign \new_Sorter100|19661_  = \new_Sorter100|19560_  | \new_Sorter100|19561_ ;
  assign \new_Sorter100|19662_  = \new_Sorter100|19562_  & \new_Sorter100|19563_ ;
  assign \new_Sorter100|19663_  = \new_Sorter100|19562_  | \new_Sorter100|19563_ ;
  assign \new_Sorter100|19664_  = \new_Sorter100|19564_  & \new_Sorter100|19565_ ;
  assign \new_Sorter100|19665_  = \new_Sorter100|19564_  | \new_Sorter100|19565_ ;
  assign \new_Sorter100|19666_  = \new_Sorter100|19566_  & \new_Sorter100|19567_ ;
  assign \new_Sorter100|19667_  = \new_Sorter100|19566_  | \new_Sorter100|19567_ ;
  assign \new_Sorter100|19668_  = \new_Sorter100|19568_  & \new_Sorter100|19569_ ;
  assign \new_Sorter100|19669_  = \new_Sorter100|19568_  | \new_Sorter100|19569_ ;
  assign \new_Sorter100|19670_  = \new_Sorter100|19570_  & \new_Sorter100|19571_ ;
  assign \new_Sorter100|19671_  = \new_Sorter100|19570_  | \new_Sorter100|19571_ ;
  assign \new_Sorter100|19672_  = \new_Sorter100|19572_  & \new_Sorter100|19573_ ;
  assign \new_Sorter100|19673_  = \new_Sorter100|19572_  | \new_Sorter100|19573_ ;
  assign \new_Sorter100|19674_  = \new_Sorter100|19574_  & \new_Sorter100|19575_ ;
  assign \new_Sorter100|19675_  = \new_Sorter100|19574_  | \new_Sorter100|19575_ ;
  assign \new_Sorter100|19676_  = \new_Sorter100|19576_  & \new_Sorter100|19577_ ;
  assign \new_Sorter100|19677_  = \new_Sorter100|19576_  | \new_Sorter100|19577_ ;
  assign \new_Sorter100|19678_  = \new_Sorter100|19578_  & \new_Sorter100|19579_ ;
  assign \new_Sorter100|19679_  = \new_Sorter100|19578_  | \new_Sorter100|19579_ ;
  assign \new_Sorter100|19680_  = \new_Sorter100|19580_  & \new_Sorter100|19581_ ;
  assign \new_Sorter100|19681_  = \new_Sorter100|19580_  | \new_Sorter100|19581_ ;
  assign \new_Sorter100|19682_  = \new_Sorter100|19582_  & \new_Sorter100|19583_ ;
  assign \new_Sorter100|19683_  = \new_Sorter100|19582_  | \new_Sorter100|19583_ ;
  assign \new_Sorter100|19684_  = \new_Sorter100|19584_  & \new_Sorter100|19585_ ;
  assign \new_Sorter100|19685_  = \new_Sorter100|19584_  | \new_Sorter100|19585_ ;
  assign \new_Sorter100|19686_  = \new_Sorter100|19586_  & \new_Sorter100|19587_ ;
  assign \new_Sorter100|19687_  = \new_Sorter100|19586_  | \new_Sorter100|19587_ ;
  assign \new_Sorter100|19688_  = \new_Sorter100|19588_  & \new_Sorter100|19589_ ;
  assign \new_Sorter100|19689_  = \new_Sorter100|19588_  | \new_Sorter100|19589_ ;
  assign \new_Sorter100|19690_  = \new_Sorter100|19590_  & \new_Sorter100|19591_ ;
  assign \new_Sorter100|19691_  = \new_Sorter100|19590_  | \new_Sorter100|19591_ ;
  assign \new_Sorter100|19692_  = \new_Sorter100|19592_  & \new_Sorter100|19593_ ;
  assign \new_Sorter100|19693_  = \new_Sorter100|19592_  | \new_Sorter100|19593_ ;
  assign \new_Sorter100|19694_  = \new_Sorter100|19594_  & \new_Sorter100|19595_ ;
  assign \new_Sorter100|19695_  = \new_Sorter100|19594_  | \new_Sorter100|19595_ ;
  assign \new_Sorter100|19696_  = \new_Sorter100|19596_  & \new_Sorter100|19597_ ;
  assign \new_Sorter100|19697_  = \new_Sorter100|19596_  | \new_Sorter100|19597_ ;
  assign \new_Sorter100|19698_  = \new_Sorter100|19598_  & \new_Sorter100|19599_ ;
  assign \new_Sorter100|19699_  = \new_Sorter100|19598_  | \new_Sorter100|19599_ ;
  assign \new_Sorter100|19700_  = \new_Sorter100|19600_ ;
  assign \new_Sorter100|19799_  = \new_Sorter100|19699_ ;
  assign \new_Sorter100|19701_  = \new_Sorter100|19601_  & \new_Sorter100|19602_ ;
  assign \new_Sorter100|19702_  = \new_Sorter100|19601_  | \new_Sorter100|19602_ ;
  assign \new_Sorter100|19703_  = \new_Sorter100|19603_  & \new_Sorter100|19604_ ;
  assign \new_Sorter100|19704_  = \new_Sorter100|19603_  | \new_Sorter100|19604_ ;
  assign \new_Sorter100|19705_  = \new_Sorter100|19605_  & \new_Sorter100|19606_ ;
  assign \new_Sorter100|19706_  = \new_Sorter100|19605_  | \new_Sorter100|19606_ ;
  assign \new_Sorter100|19707_  = \new_Sorter100|19607_  & \new_Sorter100|19608_ ;
  assign \new_Sorter100|19708_  = \new_Sorter100|19607_  | \new_Sorter100|19608_ ;
  assign \new_Sorter100|19709_  = \new_Sorter100|19609_  & \new_Sorter100|19610_ ;
  assign \new_Sorter100|19710_  = \new_Sorter100|19609_  | \new_Sorter100|19610_ ;
  assign \new_Sorter100|19711_  = \new_Sorter100|19611_  & \new_Sorter100|19612_ ;
  assign \new_Sorter100|19712_  = \new_Sorter100|19611_  | \new_Sorter100|19612_ ;
  assign \new_Sorter100|19713_  = \new_Sorter100|19613_  & \new_Sorter100|19614_ ;
  assign \new_Sorter100|19714_  = \new_Sorter100|19613_  | \new_Sorter100|19614_ ;
  assign \new_Sorter100|19715_  = \new_Sorter100|19615_  & \new_Sorter100|19616_ ;
  assign \new_Sorter100|19716_  = \new_Sorter100|19615_  | \new_Sorter100|19616_ ;
  assign \new_Sorter100|19717_  = \new_Sorter100|19617_  & \new_Sorter100|19618_ ;
  assign \new_Sorter100|19718_  = \new_Sorter100|19617_  | \new_Sorter100|19618_ ;
  assign \new_Sorter100|19719_  = \new_Sorter100|19619_  & \new_Sorter100|19620_ ;
  assign \new_Sorter100|19720_  = \new_Sorter100|19619_  | \new_Sorter100|19620_ ;
  assign \new_Sorter100|19721_  = \new_Sorter100|19621_  & \new_Sorter100|19622_ ;
  assign \new_Sorter100|19722_  = \new_Sorter100|19621_  | \new_Sorter100|19622_ ;
  assign \new_Sorter100|19723_  = \new_Sorter100|19623_  & \new_Sorter100|19624_ ;
  assign \new_Sorter100|19724_  = \new_Sorter100|19623_  | \new_Sorter100|19624_ ;
  assign \new_Sorter100|19725_  = \new_Sorter100|19625_  & \new_Sorter100|19626_ ;
  assign \new_Sorter100|19726_  = \new_Sorter100|19625_  | \new_Sorter100|19626_ ;
  assign \new_Sorter100|19727_  = \new_Sorter100|19627_  & \new_Sorter100|19628_ ;
  assign \new_Sorter100|19728_  = \new_Sorter100|19627_  | \new_Sorter100|19628_ ;
  assign \new_Sorter100|19729_  = \new_Sorter100|19629_  & \new_Sorter100|19630_ ;
  assign \new_Sorter100|19730_  = \new_Sorter100|19629_  | \new_Sorter100|19630_ ;
  assign \new_Sorter100|19731_  = \new_Sorter100|19631_  & \new_Sorter100|19632_ ;
  assign \new_Sorter100|19732_  = \new_Sorter100|19631_  | \new_Sorter100|19632_ ;
  assign \new_Sorter100|19733_  = \new_Sorter100|19633_  & \new_Sorter100|19634_ ;
  assign \new_Sorter100|19734_  = \new_Sorter100|19633_  | \new_Sorter100|19634_ ;
  assign \new_Sorter100|19735_  = \new_Sorter100|19635_  & \new_Sorter100|19636_ ;
  assign \new_Sorter100|19736_  = \new_Sorter100|19635_  | \new_Sorter100|19636_ ;
  assign \new_Sorter100|19737_  = \new_Sorter100|19637_  & \new_Sorter100|19638_ ;
  assign \new_Sorter100|19738_  = \new_Sorter100|19637_  | \new_Sorter100|19638_ ;
  assign \new_Sorter100|19739_  = \new_Sorter100|19639_  & \new_Sorter100|19640_ ;
  assign \new_Sorter100|19740_  = \new_Sorter100|19639_  | \new_Sorter100|19640_ ;
  assign \new_Sorter100|19741_  = \new_Sorter100|19641_  & \new_Sorter100|19642_ ;
  assign \new_Sorter100|19742_  = \new_Sorter100|19641_  | \new_Sorter100|19642_ ;
  assign \new_Sorter100|19743_  = \new_Sorter100|19643_  & \new_Sorter100|19644_ ;
  assign \new_Sorter100|19744_  = \new_Sorter100|19643_  | \new_Sorter100|19644_ ;
  assign \new_Sorter100|19745_  = \new_Sorter100|19645_  & \new_Sorter100|19646_ ;
  assign \new_Sorter100|19746_  = \new_Sorter100|19645_  | \new_Sorter100|19646_ ;
  assign \new_Sorter100|19747_  = \new_Sorter100|19647_  & \new_Sorter100|19648_ ;
  assign \new_Sorter100|19748_  = \new_Sorter100|19647_  | \new_Sorter100|19648_ ;
  assign \new_Sorter100|19749_  = \new_Sorter100|19649_  & \new_Sorter100|19650_ ;
  assign \new_Sorter100|19750_  = \new_Sorter100|19649_  | \new_Sorter100|19650_ ;
  assign \new_Sorter100|19751_  = \new_Sorter100|19651_  & \new_Sorter100|19652_ ;
  assign \new_Sorter100|19752_  = \new_Sorter100|19651_  | \new_Sorter100|19652_ ;
  assign \new_Sorter100|19753_  = \new_Sorter100|19653_  & \new_Sorter100|19654_ ;
  assign \new_Sorter100|19754_  = \new_Sorter100|19653_  | \new_Sorter100|19654_ ;
  assign \new_Sorter100|19755_  = \new_Sorter100|19655_  & \new_Sorter100|19656_ ;
  assign \new_Sorter100|19756_  = \new_Sorter100|19655_  | \new_Sorter100|19656_ ;
  assign \new_Sorter100|19757_  = \new_Sorter100|19657_  & \new_Sorter100|19658_ ;
  assign \new_Sorter100|19758_  = \new_Sorter100|19657_  | \new_Sorter100|19658_ ;
  assign \new_Sorter100|19759_  = \new_Sorter100|19659_  & \new_Sorter100|19660_ ;
  assign \new_Sorter100|19760_  = \new_Sorter100|19659_  | \new_Sorter100|19660_ ;
  assign \new_Sorter100|19761_  = \new_Sorter100|19661_  & \new_Sorter100|19662_ ;
  assign \new_Sorter100|19762_  = \new_Sorter100|19661_  | \new_Sorter100|19662_ ;
  assign \new_Sorter100|19763_  = \new_Sorter100|19663_  & \new_Sorter100|19664_ ;
  assign \new_Sorter100|19764_  = \new_Sorter100|19663_  | \new_Sorter100|19664_ ;
  assign \new_Sorter100|19765_  = \new_Sorter100|19665_  & \new_Sorter100|19666_ ;
  assign \new_Sorter100|19766_  = \new_Sorter100|19665_  | \new_Sorter100|19666_ ;
  assign \new_Sorter100|19767_  = \new_Sorter100|19667_  & \new_Sorter100|19668_ ;
  assign \new_Sorter100|19768_  = \new_Sorter100|19667_  | \new_Sorter100|19668_ ;
  assign \new_Sorter100|19769_  = \new_Sorter100|19669_  & \new_Sorter100|19670_ ;
  assign \new_Sorter100|19770_  = \new_Sorter100|19669_  | \new_Sorter100|19670_ ;
  assign \new_Sorter100|19771_  = \new_Sorter100|19671_  & \new_Sorter100|19672_ ;
  assign \new_Sorter100|19772_  = \new_Sorter100|19671_  | \new_Sorter100|19672_ ;
  assign \new_Sorter100|19773_  = \new_Sorter100|19673_  & \new_Sorter100|19674_ ;
  assign \new_Sorter100|19774_  = \new_Sorter100|19673_  | \new_Sorter100|19674_ ;
  assign \new_Sorter100|19775_  = \new_Sorter100|19675_  & \new_Sorter100|19676_ ;
  assign \new_Sorter100|19776_  = \new_Sorter100|19675_  | \new_Sorter100|19676_ ;
  assign \new_Sorter100|19777_  = \new_Sorter100|19677_  & \new_Sorter100|19678_ ;
  assign \new_Sorter100|19778_  = \new_Sorter100|19677_  | \new_Sorter100|19678_ ;
  assign \new_Sorter100|19779_  = \new_Sorter100|19679_  & \new_Sorter100|19680_ ;
  assign \new_Sorter100|19780_  = \new_Sorter100|19679_  | \new_Sorter100|19680_ ;
  assign \new_Sorter100|19781_  = \new_Sorter100|19681_  & \new_Sorter100|19682_ ;
  assign \new_Sorter100|19782_  = \new_Sorter100|19681_  | \new_Sorter100|19682_ ;
  assign \new_Sorter100|19783_  = \new_Sorter100|19683_  & \new_Sorter100|19684_ ;
  assign \new_Sorter100|19784_  = \new_Sorter100|19683_  | \new_Sorter100|19684_ ;
  assign \new_Sorter100|19785_  = \new_Sorter100|19685_  & \new_Sorter100|19686_ ;
  assign \new_Sorter100|19786_  = \new_Sorter100|19685_  | \new_Sorter100|19686_ ;
  assign \new_Sorter100|19787_  = \new_Sorter100|19687_  & \new_Sorter100|19688_ ;
  assign \new_Sorter100|19788_  = \new_Sorter100|19687_  | \new_Sorter100|19688_ ;
  assign \new_Sorter100|19789_  = \new_Sorter100|19689_  & \new_Sorter100|19690_ ;
  assign \new_Sorter100|19790_  = \new_Sorter100|19689_  | \new_Sorter100|19690_ ;
  assign \new_Sorter100|19791_  = \new_Sorter100|19691_  & \new_Sorter100|19692_ ;
  assign \new_Sorter100|19792_  = \new_Sorter100|19691_  | \new_Sorter100|19692_ ;
  assign \new_Sorter100|19793_  = \new_Sorter100|19693_  & \new_Sorter100|19694_ ;
  assign \new_Sorter100|19794_  = \new_Sorter100|19693_  | \new_Sorter100|19694_ ;
  assign \new_Sorter100|19795_  = \new_Sorter100|19695_  & \new_Sorter100|19696_ ;
  assign \new_Sorter100|19796_  = \new_Sorter100|19695_  | \new_Sorter100|19696_ ;
  assign \new_Sorter100|19797_  = \new_Sorter100|19697_  & \new_Sorter100|19698_ ;
  assign \new_Sorter100|19798_  = \new_Sorter100|19697_  | \new_Sorter100|19698_ ;
  assign y00 = \new_Sorter100|19700_  & \new_Sorter100|19701_ ;
  assign y01 = \new_Sorter100|19700_  | \new_Sorter100|19701_ ;
  assign y02 = \new_Sorter100|19702_  & \new_Sorter100|19703_ ;
  assign y03 = \new_Sorter100|19702_  | \new_Sorter100|19703_ ;
  assign y04 = \new_Sorter100|19704_  & \new_Sorter100|19705_ ;
  assign y05 = \new_Sorter100|19704_  | \new_Sorter100|19705_ ;
  assign y06 = \new_Sorter100|19706_  & \new_Sorter100|19707_ ;
  assign y07 = \new_Sorter100|19706_  | \new_Sorter100|19707_ ;
  assign y08 = \new_Sorter100|19708_  & \new_Sorter100|19709_ ;
  assign y09 = \new_Sorter100|19708_  | \new_Sorter100|19709_ ;
  assign y10 = \new_Sorter100|19710_  & \new_Sorter100|19711_ ;
  assign y11 = \new_Sorter100|19710_  | \new_Sorter100|19711_ ;
  assign y12 = \new_Sorter100|19712_  & \new_Sorter100|19713_ ;
  assign y13 = \new_Sorter100|19712_  | \new_Sorter100|19713_ ;
  assign y14 = \new_Sorter100|19714_  & \new_Sorter100|19715_ ;
  assign y15 = \new_Sorter100|19714_  | \new_Sorter100|19715_ ;
  assign y16 = \new_Sorter100|19716_  & \new_Sorter100|19717_ ;
  assign y17 = \new_Sorter100|19716_  | \new_Sorter100|19717_ ;
  assign y18 = \new_Sorter100|19718_  & \new_Sorter100|19719_ ;
  assign y19 = \new_Sorter100|19718_  | \new_Sorter100|19719_ ;
  assign y20 = \new_Sorter100|19720_  & \new_Sorter100|19721_ ;
  assign y21 = \new_Sorter100|19720_  | \new_Sorter100|19721_ ;
  assign y22 = \new_Sorter100|19722_  & \new_Sorter100|19723_ ;
  assign y23 = \new_Sorter100|19722_  | \new_Sorter100|19723_ ;
  assign y24 = \new_Sorter100|19724_  & \new_Sorter100|19725_ ;
  assign y25 = \new_Sorter100|19724_  | \new_Sorter100|19725_ ;
  assign y26 = \new_Sorter100|19726_  & \new_Sorter100|19727_ ;
  assign y27 = \new_Sorter100|19726_  | \new_Sorter100|19727_ ;
  assign y28 = \new_Sorter100|19728_  & \new_Sorter100|19729_ ;
  assign y29 = \new_Sorter100|19728_  | \new_Sorter100|19729_ ;
  assign y30 = \new_Sorter100|19730_  & \new_Sorter100|19731_ ;
  assign y31 = \new_Sorter100|19730_  | \new_Sorter100|19731_ ;
  assign y32 = \new_Sorter100|19732_  & \new_Sorter100|19733_ ;
  assign y33 = \new_Sorter100|19732_  | \new_Sorter100|19733_ ;
  assign y34 = \new_Sorter100|19734_  & \new_Sorter100|19735_ ;
  assign y35 = \new_Sorter100|19734_  | \new_Sorter100|19735_ ;
  assign y36 = \new_Sorter100|19736_  & \new_Sorter100|19737_ ;
  assign y37 = \new_Sorter100|19736_  | \new_Sorter100|19737_ ;
  assign y38 = \new_Sorter100|19738_  & \new_Sorter100|19739_ ;
  assign y39 = \new_Sorter100|19738_  | \new_Sorter100|19739_ ;
  assign y40 = \new_Sorter100|19740_  & \new_Sorter100|19741_ ;
  assign y41 = \new_Sorter100|19740_  | \new_Sorter100|19741_ ;
  assign y42 = \new_Sorter100|19742_  & \new_Sorter100|19743_ ;
  assign y43 = \new_Sorter100|19742_  | \new_Sorter100|19743_ ;
  assign y44 = \new_Sorter100|19744_  & \new_Sorter100|19745_ ;
  assign y45 = \new_Sorter100|19744_  | \new_Sorter100|19745_ ;
  assign y46 = \new_Sorter100|19746_  & \new_Sorter100|19747_ ;
  assign y47 = \new_Sorter100|19746_  | \new_Sorter100|19747_ ;
  assign y48 = \new_Sorter100|19748_  & \new_Sorter100|19749_ ;
  assign y49 = \new_Sorter100|19748_  | \new_Sorter100|19749_ ;
  assign y50 = \new_Sorter100|19750_  & \new_Sorter100|19751_ ;
  assign y51 = \new_Sorter100|19750_  | \new_Sorter100|19751_ ;
  assign y52 = \new_Sorter100|19752_  & \new_Sorter100|19753_ ;
  assign y53 = \new_Sorter100|19752_  | \new_Sorter100|19753_ ;
  assign y54 = \new_Sorter100|19754_  & \new_Sorter100|19755_ ;
  assign y55 = \new_Sorter100|19754_  | \new_Sorter100|19755_ ;
  assign y56 = \new_Sorter100|19756_  & \new_Sorter100|19757_ ;
  assign y57 = \new_Sorter100|19756_  | \new_Sorter100|19757_ ;
  assign y58 = \new_Sorter100|19758_  & \new_Sorter100|19759_ ;
  assign y59 = \new_Sorter100|19758_  | \new_Sorter100|19759_ ;
  assign y60 = \new_Sorter100|19760_  & \new_Sorter100|19761_ ;
  assign y61 = \new_Sorter100|19760_  | \new_Sorter100|19761_ ;
  assign y62 = \new_Sorter100|19762_  & \new_Sorter100|19763_ ;
  assign y63 = \new_Sorter100|19762_  | \new_Sorter100|19763_ ;
  assign y64 = \new_Sorter100|19764_  & \new_Sorter100|19765_ ;
  assign y65 = \new_Sorter100|19764_  | \new_Sorter100|19765_ ;
  assign y66 = \new_Sorter100|19766_  & \new_Sorter100|19767_ ;
  assign y67 = \new_Sorter100|19766_  | \new_Sorter100|19767_ ;
  assign y68 = \new_Sorter100|19768_  & \new_Sorter100|19769_ ;
  assign y69 = \new_Sorter100|19768_  | \new_Sorter100|19769_ ;
  assign y70 = \new_Sorter100|19770_  & \new_Sorter100|19771_ ;
  assign y71 = \new_Sorter100|19770_  | \new_Sorter100|19771_ ;
  assign y72 = \new_Sorter100|19772_  & \new_Sorter100|19773_ ;
  assign y73 = \new_Sorter100|19772_  | \new_Sorter100|19773_ ;
  assign y74 = \new_Sorter100|19774_  & \new_Sorter100|19775_ ;
  assign y75 = \new_Sorter100|19774_  | \new_Sorter100|19775_ ;
  assign y76 = \new_Sorter100|19776_  & \new_Sorter100|19777_ ;
  assign y77 = \new_Sorter100|19776_  | \new_Sorter100|19777_ ;
  assign y78 = \new_Sorter100|19778_  & \new_Sorter100|19779_ ;
  assign y79 = \new_Sorter100|19778_  | \new_Sorter100|19779_ ;
  assign y80 = \new_Sorter100|19780_  & \new_Sorter100|19781_ ;
  assign y81 = \new_Sorter100|19780_  | \new_Sorter100|19781_ ;
  assign y82 = \new_Sorter100|19782_  & \new_Sorter100|19783_ ;
  assign y83 = \new_Sorter100|19782_  | \new_Sorter100|19783_ ;
  assign y84 = \new_Sorter100|19784_  & \new_Sorter100|19785_ ;
  assign y85 = \new_Sorter100|19784_  | \new_Sorter100|19785_ ;
  assign y86 = \new_Sorter100|19786_  & \new_Sorter100|19787_ ;
  assign y87 = \new_Sorter100|19786_  | \new_Sorter100|19787_ ;
  assign y88 = \new_Sorter100|19788_  & \new_Sorter100|19789_ ;
  assign y89 = \new_Sorter100|19788_  | \new_Sorter100|19789_ ;
  assign y90 = \new_Sorter100|19790_  & \new_Sorter100|19791_ ;
  assign y91 = \new_Sorter100|19790_  | \new_Sorter100|19791_ ;
  assign y92 = \new_Sorter100|19792_  & \new_Sorter100|19793_ ;
  assign y93 = \new_Sorter100|19792_  | \new_Sorter100|19793_ ;
  assign y94 = \new_Sorter100|19794_  & \new_Sorter100|19795_ ;
  assign y95 = \new_Sorter100|19794_  | \new_Sorter100|19795_ ;
  assign y96 = \new_Sorter100|19796_  & \new_Sorter100|19797_ ;
  assign y97 = \new_Sorter100|19796_  | \new_Sorter100|19797_ ;
  assign y98 = \new_Sorter100|19798_  & \new_Sorter100|19799_ ;
  assign y99 = \new_Sorter100|19798_  | \new_Sorter100|19799_ ;
endmodule


