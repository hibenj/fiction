// Benchmark "Multi8" written by ABC on Tue Apr  9 09:18:12 2024

module Multi8 ( 
    a0, a1, a2, a3, a4, a5, a6, a7, b0, b1, b2, b3, b4, b5, b6, b7,
    m00, m01, m02, m03, m04, m05, m06, m07, m08, m09, m10, m11, m12, m13,
    m14, m15  );
  input  a0, a1, a2, a3, a4, a5, a6, a7, b0, b1, b2, b3, b4, b5, b6, b7;
  output m00, m01, m02, m03, m04, m05, m06, m07, m08, m09, m10, m11, m12, m13,
    m14, m15;
  wire new_n246_, new_n248_, new_n250_, new_n252_, new_n254_, new_n256_,
    new_n258_, new_n260_, new_n262_, new_n264_, new_n266_, new_n268_,
    new_n270_, new_n272_, new_n274_, new_n276_, new_n278_, new_n280_,
    new_n282_, new_n284_, new_n286_, new_n288_, new_n290_, new_n292_,
    new_n294_, new_n296_, new_n298_, new_n300_, new_n302_, new_n304_,
    new_n306_, new_n308_, new_n310_, new_n312_, new_n314_, new_n316_,
    new_n318_, new_n320_, new_n322_, new_n324_, new_n326_, new_n328_,
    new_n330_, new_n332_, new_n334_, new_n336_, new_n338_, new_n340_,
    new_n342_, new_n344_, new_n346_, new_n348_, new_n350_, new_n352_,
    new_n354_, new_n356_, new_n358_, new_n360_, new_n362_, new_n364_,
    new_n366_, new_n368_, new_n370_, new_n372_, new_n374_, new_n376_,
    new_n378_, new_n380_, new_n382_, new_n384_, new_n386_, new_n388_,
    new_n390_, new_n392_, new_n394_, new_n396_, new_n398_, new_n400_,
    new_n402_, new_n404_, new_n406_, new_n408_, new_n410_, new_n412_,
    new_n414_, new_n416_, new_n418_, new_n420_, new_n422_, new_n424_,
    new_n426_, new_n428_, new_n430_, new_n432_, new_n434_, new_n436_,
    new_n438_, new_n440_, new_n442_, new_n444_, new_n446_, new_n448_,
    new_n450_, new_n452_, new_n454_, new_n456_, new_n458_, new_n460_,
    new_n462_, new_n464_, new_n466_, new_n468_, new_n470_, new_n472_,
    new_n474_, new_n476_, new_n478_, new_n480_, new_n482_, new_n484_,
    new_n486_, new_n488_, new_n490_, new_n492_, new_n494_, new_n496_,
    new_n498_, new_n500_, new_n502_, new_n504_, new_n506_, new_n508_,
    new_n510_, new_n512_, new_n514_, new_n516_, new_n518_, new_n520_,
    new_n522_, new_n524_, new_n526_, new_n528_, new_n530_, new_n532_,
    new_n534_, new_n536_, new_n538_, new_n540_, new_n542_, new_n544_,
    new_n546_, new_n548_, new_n550_, new_n552_, new_n554_, new_n556_,
    new_n558_, new_n560_, new_n562_, new_n564_, new_n566_, new_n568_,
    new_n570_, new_n572_, new_n574_, new_n576_, new_n578_, new_n580_,
    new_n582_, new_n584_, new_n586_, new_n588_, new_n590_, new_n592_,
    new_n594_, new_n596_, new_n598_, new_n600_, new_n602_, new_n604_,
    new_n606_, new_n608_, new_n610_, new_n612_, new_n614_, new_n616_,
    new_n618_, new_n620_, new_n622_, new_n624_, new_n626_, new_n628_,
    new_n630_, new_n632_, new_n634_, new_n636_, new_n638_, new_n640_,
    new_n642_, new_n644_, new_n646_, new_n648_, new_n650_, new_n652_,
    new_n654_, new_n656_, new_n658_, new_n660_, new_n662_, new_n664_,
    new_n666_, new_n668_, new_n670_, new_n672_, new_n674_, new_n676_,
    new_n678_, new_n680_, new_n682_, new_n684_, new_n686_, new_n688_,
    new_n690_, new_n692_, new_n694_, new_n696_, new_n698_, new_n700_,
    new_n702_, new_n704_, new_n706_, new_n708_, new_n710_, new_n712_,
    new_n714_, new_n716_, new_n718_, new_n720_, new_n722_, new_n724_,
    new_n726_, new_n728_, new_n730_, new_n732_, new_n734_, new_n736_,
    new_n738_, new_n740_, new_n742_, new_n744_, new_n746_, new_n748_,
    new_n750_, new_n752_, new_n754_, new_n756_, new_n758_, new_n760_,
    new_n762_, new_n764_, new_n766_, new_n768_, new_n770_, new_n772_,
    new_n774_, new_n776_, new_n778_, new_n780_, new_n782_, new_n784_,
    new_n786_, new_n788_, new_n790_, new_n792_, new_n794_, new_n796_,
    new_n798_, new_n800_, new_n802_, new_n804_, new_n806_, new_n808_,
    new_n810_, new_n812_, new_n814_, new_n816_, new_n818_, new_n820_,
    new_n822_, new_n824_, new_n826_, new_n828_, new_n830_, new_n832_,
    new_n834_, new_n836_, new_n838_, new_n840_, new_n842_, new_n844_,
    new_n846_, new_n848_, new_n850_, new_n852_, new_n854_, new_n856_,
    new_n858_, new_n860_, new_n862_, new_n864_, new_n866_, new_n868_,
    new_n870_, new_n872_, new_n874_, new_n876_, new_n878_, new_n880_,
    new_n882_, new_n884_, new_n886_, new_n888_, new_n890_, new_n892_,
    new_n894_, new_n896_, new_n898_, new_n900_, new_n902_, new_n904_,
    new_n906_, new_n908_, new_n910_, new_n912_, new_n914_, new_n916_,
    new_n918_, new_n920_, new_n922_, new_n924_, new_n926_, new_n928_,
    new_n930_, new_n932_, new_n934_, new_n936_, new_n938_, new_n940_,
    new_n942_, new_n944_, \new_Multi8|y0_00_ , \new_Multi8|y0_01_ ,
    \new_Multi8|y0_02_ , \new_Multi8|y0_03_ , \new_Multi8|y0_04_ ,
    \new_Multi8|y0_05_ , \new_Multi8|y0_06_ , \new_Multi8|y0_07_ ,
    \new_Multi8|y0_08_ , \new_Multi8|y0_09_ , \new_Multi8|y0_10_ ,
    \new_Multi8|y0_11_ , \new_Multi8|y0_12_ , \new_Multi8|y0_13_ ,
    \new_Multi8|y0_14_ , \new_Multi8|y0_15_ , \new_Multi8|y1_00_ ,
    \new_Multi8|y1_01_ , \new_Multi8|y1_02_ , \new_Multi8|y1_03_ ,
    \new_Multi8|y1_04_ , \new_Multi8|y1_05_ , \new_Multi8|y1_06_ ,
    \new_Multi8|y1_07_ , \new_Multi8|y1_08_ , \new_Multi8|y1_09_ ,
    \new_Multi8|y1_10_ , \new_Multi8|y1_11_ , \new_Multi8|y1_12_ ,
    \new_Multi8|y1_13_ , \new_Multi8|y1_14_ , \new_Multi8|y1_15_ ,
    \new_Multi8|y2_00_ , \new_Multi8|y2_01_ , \new_Multi8|y2_02_ ,
    \new_Multi8|y2_03_ , \new_Multi8|y2_04_ , \new_Multi8|y2_05_ ,
    \new_Multi8|y2_06_ , \new_Multi8|y2_07_ , \new_Multi8|y2_08_ ,
    \new_Multi8|y2_09_ , \new_Multi8|y2_10_ , \new_Multi8|y2_11_ ,
    \new_Multi8|y2_12_ , \new_Multi8|y2_13_ , \new_Multi8|y2_14_ ,
    \new_Multi8|y2_15_ , \new_Multi8|y3_00_ , \new_Multi8|y3_01_ ,
    \new_Multi8|y3_02_ , \new_Multi8|y3_03_ , \new_Multi8|y3_04_ ,
    \new_Multi8|y3_05_ , \new_Multi8|y3_06_ , \new_Multi8|y3_07_ ,
    \new_Multi8|y3_08_ , \new_Multi8|y3_09_ , \new_Multi8|y3_10_ ,
    \new_Multi8|y3_11_ , \new_Multi8|y3_12_ , \new_Multi8|y3_13_ ,
    \new_Multi8|y3_14_ , \new_Multi8|y3_15_ , \new_Multi8|y4_00_ ,
    \new_Multi8|y4_01_ , \new_Multi8|y4_02_ , \new_Multi8|y4_03_ ,
    \new_Multi8|y4_04_ , \new_Multi8|y4_05_ , \new_Multi8|y4_06_ ,
    \new_Multi8|y4_07_ , \new_Multi8|y4_08_ , \new_Multi8|y4_09_ ,
    \new_Multi8|y4_10_ , \new_Multi8|y4_11_ , \new_Multi8|y4_12_ ,
    \new_Multi8|y4_13_ , \new_Multi8|y4_14_ , \new_Multi8|y4_15_ ,
    \new_Multi8|x0_00_ , \new_Multi8|x0_01_ , \new_Multi8|x0_02_ ,
    \new_Multi8|x0_03_ , \new_Multi8|x0_04_ , \new_Multi8|x0_05_ ,
    \new_Multi8|x0_06_ , \new_Multi8|x0_07_ , \new_Multi8|x0_08_ ,
    \new_Multi8|x0_09_ , \new_Multi8|x0_10_ , \new_Multi8|x0_11_ ,
    \new_Multi8|x0_12_ , \new_Multi8|x0_13_ , \new_Multi8|x0_14_ ,
    \new_Multi8|x0_15_ , \new_Multi8|ADD16(1)|c_ , new_n1075_, new_n1077_,
    new_n1079_, new_n1081_, new_n1083_, \new_Multi8|x1_00_ ,
    \new_Multi8|ADD16(1)|00_ , new_n1087_, new_n1089_, new_n1091_,
    new_n1093_, new_n1095_, \new_Multi8|x1_01_ , \new_Multi8|ADD16(1)|01_ ,
    new_n1099_, new_n1101_, new_n1103_, new_n1105_, new_n1107_,
    \new_Multi8|x1_02_ , \new_Multi8|ADD16(1)|02_ , new_n1111_, new_n1113_,
    new_n1115_, new_n1117_, new_n1119_, \new_Multi8|x1_03_ ,
    \new_Multi8|ADD16(1)|03_ , new_n1123_, new_n1125_, new_n1127_,
    new_n1129_, new_n1131_, \new_Multi8|x1_04_ , \new_Multi8|ADD16(1)|04_ ,
    new_n1135_, new_n1137_, new_n1139_, new_n1141_, new_n1143_,
    \new_Multi8|x1_05_ , \new_Multi8|ADD16(1)|05_ , new_n1147_, new_n1149_,
    new_n1151_, new_n1153_, new_n1155_, \new_Multi8|x1_06_ ,
    \new_Multi8|ADD16(1)|06_ , new_n1159_, new_n1161_, new_n1163_,
    new_n1165_, new_n1167_, \new_Multi8|x1_07_ , \new_Multi8|ADD16(1)|07_ ,
    new_n1171_, new_n1173_, new_n1175_, new_n1177_, new_n1179_,
    \new_Multi8|x1_08_ , \new_Multi8|ADD16(1)|08_ , new_n1183_, new_n1185_,
    new_n1187_, new_n1189_, new_n1191_, \new_Multi8|x1_09_ ,
    \new_Multi8|ADD16(1)|09_ , new_n1195_, new_n1197_, new_n1199_,
    new_n1201_, new_n1203_, \new_Multi8|x1_10_ , \new_Multi8|ADD16(1)|10_ ,
    new_n1207_, new_n1209_, new_n1211_, new_n1213_, new_n1215_,
    \new_Multi8|x1_11_ , \new_Multi8|ADD16(1)|11_ , new_n1219_, new_n1221_,
    new_n1223_, new_n1225_, new_n1227_, \new_Multi8|x1_12_ ,
    \new_Multi8|ADD16(1)|12_ , new_n1231_, new_n1233_, new_n1235_,
    new_n1237_, new_n1239_, \new_Multi8|x1_13_ , \new_Multi8|ADD16(1)|13_ ,
    new_n1243_, new_n1245_, new_n1247_, new_n1249_, new_n1251_,
    \new_Multi8|x1_14_ , \new_Multi8|ADD16(1)|14_ , new_n1255_, new_n1257_,
    new_n1259_, new_n1261_, new_n1263_, \new_Multi8|x1_15_ ,
    \new_Multi8|ADD16(18)|c_ , new_n1284_, new_n1286_, new_n1288_,
    new_n1290_, new_n1292_, \new_Multi8|x2_00_ ,
    \new_Multi8|ADD16(18)|00_ , new_n1296_, new_n1298_, new_n1300_,
    new_n1302_, new_n1304_, \new_Multi8|x2_01_ ,
    \new_Multi8|ADD16(18)|01_ , new_n1308_, new_n1310_, new_n1312_,
    new_n1314_, new_n1316_, \new_Multi8|x2_02_ ,
    \new_Multi8|ADD16(18)|02_ , new_n1320_, new_n1322_, new_n1324_,
    new_n1326_, new_n1328_, \new_Multi8|x2_03_ ,
    \new_Multi8|ADD16(18)|03_ , new_n1332_, new_n1334_, new_n1336_,
    new_n1338_, new_n1340_, \new_Multi8|x2_04_ ,
    \new_Multi8|ADD16(18)|04_ , new_n1344_, new_n1346_, new_n1348_,
    new_n1350_, new_n1352_, \new_Multi8|x2_05_ ,
    \new_Multi8|ADD16(18)|05_ , new_n1356_, new_n1358_, new_n1360_,
    new_n1362_, new_n1364_, \new_Multi8|x2_06_ ,
    \new_Multi8|ADD16(18)|06_ , new_n1368_, new_n1370_, new_n1372_,
    new_n1374_, new_n1376_, \new_Multi8|x2_07_ ,
    \new_Multi8|ADD16(18)|07_ , new_n1380_, new_n1382_, new_n1384_,
    new_n1386_, new_n1388_, \new_Multi8|x2_08_ ,
    \new_Multi8|ADD16(18)|08_ , new_n1392_, new_n1394_, new_n1396_,
    new_n1398_, new_n1400_, \new_Multi8|x2_09_ ,
    \new_Multi8|ADD16(18)|09_ , new_n1404_, new_n1406_, new_n1408_,
    new_n1410_, new_n1412_, \new_Multi8|x2_10_ ,
    \new_Multi8|ADD16(18)|10_ , new_n1416_, new_n1418_, new_n1420_,
    new_n1422_, new_n1424_, \new_Multi8|x2_11_ ,
    \new_Multi8|ADD16(18)|11_ , new_n1428_, new_n1430_, new_n1432_,
    new_n1434_, new_n1436_, \new_Multi8|x2_12_ ,
    \new_Multi8|ADD16(18)|12_ , new_n1440_, new_n1442_, new_n1444_,
    new_n1446_, new_n1448_, \new_Multi8|x2_13_ ,
    \new_Multi8|ADD16(18)|13_ , new_n1452_, new_n1454_, new_n1456_,
    new_n1458_, new_n1460_, \new_Multi8|x2_14_ ,
    \new_Multi8|ADD16(18)|14_ , new_n1464_, new_n1466_, new_n1468_,
    new_n1470_, new_n1472_, \new_Multi8|x2_15_ , \new_Multi8|ADD16(35)|c_ ,
    new_n1493_, new_n1495_, new_n1497_, new_n1499_, new_n1501_,
    \new_Multi8|x3_00_ , \new_Multi8|ADD16(35)|00_ , new_n1505_,
    new_n1507_, new_n1509_, new_n1511_, new_n1513_, \new_Multi8|x3_01_ ,
    \new_Multi8|ADD16(35)|01_ , new_n1517_, new_n1519_, new_n1521_,
    new_n1523_, new_n1525_, \new_Multi8|x3_02_ ,
    \new_Multi8|ADD16(35)|02_ , new_n1529_, new_n1531_, new_n1533_,
    new_n1535_, new_n1537_, \new_Multi8|x3_03_ ,
    \new_Multi8|ADD16(35)|03_ , new_n1541_, new_n1543_, new_n1545_,
    new_n1547_, new_n1549_, \new_Multi8|x3_04_ ,
    \new_Multi8|ADD16(35)|04_ , new_n1553_, new_n1555_, new_n1557_,
    new_n1559_, new_n1561_, \new_Multi8|x3_05_ ,
    \new_Multi8|ADD16(35)|05_ , new_n1565_, new_n1567_, new_n1569_,
    new_n1571_, new_n1573_, \new_Multi8|x3_06_ ,
    \new_Multi8|ADD16(35)|06_ , new_n1577_, new_n1579_, new_n1581_,
    new_n1583_, new_n1585_, \new_Multi8|x3_07_ ,
    \new_Multi8|ADD16(35)|07_ , new_n1589_, new_n1591_, new_n1593_,
    new_n1595_, new_n1597_, \new_Multi8|x3_08_ ,
    \new_Multi8|ADD16(35)|08_ , new_n1601_, new_n1603_, new_n1605_,
    new_n1607_, new_n1609_, \new_Multi8|x3_09_ ,
    \new_Multi8|ADD16(35)|09_ , new_n1613_, new_n1615_, new_n1617_,
    new_n1619_, new_n1621_, \new_Multi8|x3_10_ ,
    \new_Multi8|ADD16(35)|10_ , new_n1625_, new_n1627_, new_n1629_,
    new_n1631_, new_n1633_, \new_Multi8|x3_11_ ,
    \new_Multi8|ADD16(35)|11_ , new_n1637_, new_n1639_, new_n1641_,
    new_n1643_, new_n1645_, \new_Multi8|x3_12_ ,
    \new_Multi8|ADD16(35)|12_ , new_n1649_, new_n1651_, new_n1653_,
    new_n1655_, new_n1657_, \new_Multi8|x3_13_ ,
    \new_Multi8|ADD16(35)|13_ , new_n1661_, new_n1663_, new_n1665_,
    new_n1667_, new_n1669_, \new_Multi8|x3_14_ ,
    \new_Multi8|ADD16(35)|14_ , new_n1673_, new_n1675_, new_n1677_,
    new_n1679_, new_n1681_, \new_Multi8|x3_15_ , \new_Multi8|ADD16(52)|c_ ,
    new_n1702_, new_n1704_, new_n1706_, new_n1708_, new_n1710_,
    \new_Multi8|x4_00_ , \new_Multi8|ADD16(52)|00_ , new_n1714_,
    new_n1716_, new_n1718_, new_n1720_, new_n1722_, \new_Multi8|x4_01_ ,
    \new_Multi8|ADD16(52)|01_ , new_n1726_, new_n1728_, new_n1730_,
    new_n1732_, new_n1734_, \new_Multi8|x4_02_ ,
    \new_Multi8|ADD16(52)|02_ , new_n1738_, new_n1740_, new_n1742_,
    new_n1744_, new_n1746_, \new_Multi8|x4_03_ ,
    \new_Multi8|ADD16(52)|03_ , new_n1750_, new_n1752_, new_n1754_,
    new_n1756_, new_n1758_, \new_Multi8|x4_04_ ,
    \new_Multi8|ADD16(52)|04_ , new_n1762_, new_n1764_, new_n1766_,
    new_n1768_, new_n1770_, \new_Multi8|x4_05_ ,
    \new_Multi8|ADD16(52)|05_ , new_n1774_, new_n1776_, new_n1778_,
    new_n1780_, new_n1782_, \new_Multi8|x4_06_ ,
    \new_Multi8|ADD16(52)|06_ , new_n1786_, new_n1788_, new_n1790_,
    new_n1792_, new_n1794_, \new_Multi8|x4_07_ ,
    \new_Multi8|ADD16(52)|07_ , new_n1798_, new_n1800_, new_n1802_,
    new_n1804_, new_n1806_, \new_Multi8|x4_08_ ,
    \new_Multi8|ADD16(52)|08_ , new_n1810_, new_n1812_, new_n1814_,
    new_n1816_, new_n1818_, \new_Multi8|x4_09_ ,
    \new_Multi8|ADD16(52)|09_ , new_n1822_, new_n1824_, new_n1826_,
    new_n1828_, new_n1830_, \new_Multi8|x4_10_ ,
    \new_Multi8|ADD16(52)|10_ , new_n1834_, new_n1836_, new_n1838_,
    new_n1840_, new_n1842_, \new_Multi8|x4_11_ ,
    \new_Multi8|ADD16(52)|11_ , new_n1846_, new_n1848_, new_n1850_,
    new_n1852_, new_n1854_, \new_Multi8|x4_12_ ,
    \new_Multi8|ADD16(52)|12_ , new_n1858_, new_n1860_, new_n1862_,
    new_n1864_, new_n1866_, \new_Multi8|x4_13_ ,
    \new_Multi8|ADD16(52)|13_ , new_n1870_, new_n1872_, new_n1874_,
    new_n1876_, new_n1878_, \new_Multi8|x4_14_ ,
    \new_Multi8|ADD16(52)|14_ , new_n1882_, new_n1884_, new_n1886_,
    new_n1888_, new_n1890_, \new_Multi8|x4_15_ , \new_Multi8|ADD16(69)|c_ ,
    new_n1911_, new_n1913_, new_n1915_, new_n1917_, new_n1919_,
    \new_Multi8|x5_00_ , \new_Multi8|ADD16(69)|00_ , new_n1923_,
    new_n1925_, new_n1927_, new_n1929_, new_n1931_, \new_Multi8|x5_01_ ,
    \new_Multi8|ADD16(69)|01_ , new_n1935_, new_n1937_, new_n1939_,
    new_n1941_, new_n1943_, \new_Multi8|x5_02_ ,
    \new_Multi8|ADD16(69)|02_ , new_n1947_, new_n1949_, new_n1951_,
    new_n1953_, new_n1955_, \new_Multi8|x5_03_ ,
    \new_Multi8|ADD16(69)|03_ , new_n1959_, new_n1961_, new_n1963_,
    new_n1965_, new_n1967_, \new_Multi8|x5_04_ ,
    \new_Multi8|ADD16(69)|04_ , new_n1971_, new_n1973_, new_n1975_,
    new_n1977_, new_n1979_, \new_Multi8|x5_05_ ,
    \new_Multi8|ADD16(69)|05_ , new_n1983_, new_n1985_, new_n1987_,
    new_n1989_, new_n1991_, \new_Multi8|x5_06_ ,
    \new_Multi8|ADD16(69)|06_ , new_n1995_, new_n1997_, new_n1999_,
    new_n2001_, new_n2003_, \new_Multi8|x5_07_ ,
    \new_Multi8|ADD16(69)|07_ , new_n2007_, new_n2009_, new_n2011_,
    new_n2013_, new_n2015_, \new_Multi8|x5_08_ ,
    \new_Multi8|ADD16(69)|08_ , new_n2019_, new_n2021_, new_n2023_,
    new_n2025_, new_n2027_, \new_Multi8|x5_09_ ,
    \new_Multi8|ADD16(69)|09_ , new_n2031_, new_n2033_, new_n2035_,
    new_n2037_, new_n2039_, \new_Multi8|x5_10_ ,
    \new_Multi8|ADD16(69)|10_ , new_n2043_, new_n2045_, new_n2047_,
    new_n2049_, new_n2051_, \new_Multi8|x5_11_ ,
    \new_Multi8|ADD16(69)|11_ , new_n2055_, new_n2057_, new_n2059_,
    new_n2061_, new_n2063_, \new_Multi8|x5_12_ ,
    \new_Multi8|ADD16(69)|12_ , new_n2067_, new_n2069_, new_n2071_,
    new_n2073_, new_n2075_, \new_Multi8|x5_13_ ,
    \new_Multi8|ADD16(69)|13_ , new_n2079_, new_n2081_, new_n2083_,
    new_n2085_, new_n2087_, \new_Multi8|x5_14_ ,
    \new_Multi8|ADD16(69)|14_ , new_n2091_, new_n2093_, new_n2095_,
    new_n2097_, new_n2099_, \new_Multi8|x5_15_ ;
  assign new_n246_ = 1'b0;
  assign new_n248_ = a0;
  assign new_n250_ = a1;
  assign new_n252_ = a2;
  assign new_n254_ = a3;
  assign new_n256_ = a4;
  assign new_n258_ = a5;
  assign new_n260_ = a6;
  assign new_n262_ = a7;
  assign new_n264_ = b0;
  assign new_n266_ = b1;
  assign new_n268_ = b2;
  assign new_n270_ = b3;
  assign new_n272_ = b4;
  assign new_n274_ = b5;
  assign new_n276_ = b6;
  assign new_n278_ = b7;
  assign new_n280_ = new_n264_ & ~new_n266_;
  assign new_n282_ = ~new_n264_ & new_n266_;
  assign new_n284_ = ~new_n280_ & ~new_n282_;
  assign new_n286_ = new_n248_ & new_n264_;
  assign new_n288_ = ~new_n284_ & new_n286_;
  assign new_n290_ = new_n284_ & ~new_n286_;
  assign new_n292_ = ~new_n288_ & ~new_n290_;
  assign new_n294_ = new_n264_ & ~new_n292_;
  assign new_n296_ = ~new_n264_ & new_n292_;
  assign new_n298_ = ~new_n294_ & ~new_n296_;
  assign new_n300_ = new_n248_ & ~new_n264_;
  assign new_n302_ = new_n250_ & new_n264_;
  assign new_n304_ = ~new_n284_ & ~new_n300_;
  assign new_n306_ = new_n302_ & ~new_n304_;
  assign new_n308_ = ~new_n302_ & new_n304_;
  assign new_n310_ = ~new_n306_ & ~new_n308_;
  assign new_n312_ = new_n264_ & ~new_n310_;
  assign new_n314_ = ~new_n264_ & new_n310_;
  assign new_n316_ = ~new_n312_ & ~new_n314_;
  assign new_n318_ = new_n250_ & ~new_n264_;
  assign new_n320_ = new_n252_ & new_n264_;
  assign new_n322_ = ~new_n284_ & ~new_n318_;
  assign new_n324_ = new_n320_ & ~new_n322_;
  assign new_n326_ = ~new_n320_ & new_n322_;
  assign new_n328_ = ~new_n324_ & ~new_n326_;
  assign new_n330_ = new_n264_ & ~new_n328_;
  assign new_n332_ = ~new_n264_ & new_n328_;
  assign new_n334_ = ~new_n330_ & ~new_n332_;
  assign new_n336_ = new_n252_ & ~new_n264_;
  assign new_n338_ = new_n254_ & new_n264_;
  assign new_n340_ = ~new_n284_ & ~new_n336_;
  assign new_n342_ = new_n338_ & ~new_n340_;
  assign new_n344_ = ~new_n338_ & new_n340_;
  assign new_n346_ = ~new_n342_ & ~new_n344_;
  assign new_n348_ = new_n264_ & ~new_n346_;
  assign new_n350_ = ~new_n264_ & new_n346_;
  assign new_n352_ = ~new_n348_ & ~new_n350_;
  assign new_n354_ = new_n254_ & ~new_n264_;
  assign new_n356_ = new_n256_ & new_n264_;
  assign new_n358_ = ~new_n284_ & ~new_n354_;
  assign new_n360_ = new_n356_ & ~new_n358_;
  assign new_n362_ = ~new_n356_ & new_n358_;
  assign new_n364_ = ~new_n360_ & ~new_n362_;
  assign new_n366_ = new_n264_ & ~new_n364_;
  assign new_n368_ = ~new_n264_ & new_n364_;
  assign new_n370_ = ~new_n366_ & ~new_n368_;
  assign new_n372_ = new_n256_ & ~new_n264_;
  assign new_n374_ = new_n258_ & new_n264_;
  assign new_n376_ = ~new_n284_ & ~new_n372_;
  assign new_n378_ = new_n374_ & ~new_n376_;
  assign new_n380_ = ~new_n374_ & new_n376_;
  assign new_n382_ = ~new_n378_ & ~new_n380_;
  assign new_n384_ = new_n264_ & ~new_n382_;
  assign new_n386_ = ~new_n264_ & new_n382_;
  assign new_n388_ = ~new_n384_ & ~new_n386_;
  assign new_n390_ = new_n258_ & ~new_n264_;
  assign new_n392_ = new_n260_ & new_n264_;
  assign new_n394_ = ~new_n284_ & ~new_n390_;
  assign new_n396_ = new_n392_ & ~new_n394_;
  assign new_n398_ = ~new_n392_ & new_n394_;
  assign new_n400_ = ~new_n396_ & ~new_n398_;
  assign new_n402_ = new_n264_ & ~new_n400_;
  assign new_n404_ = ~new_n264_ & new_n400_;
  assign new_n406_ = ~new_n402_ & ~new_n404_;
  assign new_n408_ = new_n260_ & ~new_n264_;
  assign new_n410_ = new_n262_ & new_n264_;
  assign new_n412_ = ~new_n284_ & ~new_n408_;
  assign new_n414_ = new_n410_ & ~new_n412_;
  assign new_n416_ = ~new_n410_ & new_n412_;
  assign new_n418_ = ~new_n414_ & ~new_n416_;
  assign new_n420_ = new_n264_ & ~new_n418_;
  assign new_n422_ = ~new_n264_ & new_n418_;
  assign new_n424_ = ~new_n420_ & ~new_n422_;
  assign new_n426_ = new_n262_ & ~new_n264_;
  assign new_n428_ = ~new_n284_ & ~new_n426_;
  assign new_n430_ = new_n410_ & ~new_n428_;
  assign new_n432_ = ~new_n410_ & new_n428_;
  assign new_n434_ = ~new_n430_ & ~new_n432_;
  assign new_n436_ = new_n264_ & ~new_n434_;
  assign new_n438_ = ~new_n264_ & new_n434_;
  assign new_n440_ = ~new_n436_ & ~new_n438_;
  assign new_n442_ = new_n268_ & ~new_n270_;
  assign new_n444_ = ~new_n268_ & new_n270_;
  assign new_n446_ = ~new_n442_ & ~new_n444_;
  assign new_n448_ = new_n266_ & ~new_n268_;
  assign new_n450_ = ~new_n266_ & new_n268_;
  assign new_n452_ = ~new_n448_ & ~new_n450_;
  assign new_n454_ = new_n248_ & ~new_n452_;
  assign new_n456_ = ~new_n446_ & new_n454_;
  assign new_n458_ = new_n446_ & ~new_n454_;
  assign new_n460_ = ~new_n456_ & ~new_n458_;
  assign new_n462_ = new_n268_ & ~new_n460_;
  assign new_n464_ = ~new_n268_ & new_n460_;
  assign new_n466_ = ~new_n462_ & ~new_n464_;
  assign new_n468_ = new_n248_ & new_n452_;
  assign new_n470_ = new_n250_ & ~new_n452_;
  assign new_n472_ = ~new_n446_ & ~new_n468_;
  assign new_n474_ = new_n470_ & ~new_n472_;
  assign new_n476_ = ~new_n470_ & new_n472_;
  assign new_n478_ = ~new_n474_ & ~new_n476_;
  assign new_n480_ = new_n268_ & ~new_n478_;
  assign new_n482_ = ~new_n268_ & new_n478_;
  assign new_n484_ = ~new_n480_ & ~new_n482_;
  assign new_n486_ = new_n250_ & new_n452_;
  assign new_n488_ = new_n252_ & ~new_n452_;
  assign new_n490_ = ~new_n446_ & ~new_n486_;
  assign new_n492_ = new_n488_ & ~new_n490_;
  assign new_n494_ = ~new_n488_ & new_n490_;
  assign new_n496_ = ~new_n492_ & ~new_n494_;
  assign new_n498_ = new_n268_ & ~new_n496_;
  assign new_n500_ = ~new_n268_ & new_n496_;
  assign new_n502_ = ~new_n498_ & ~new_n500_;
  assign new_n504_ = new_n252_ & new_n452_;
  assign new_n506_ = new_n254_ & ~new_n452_;
  assign new_n508_ = ~new_n446_ & ~new_n504_;
  assign new_n510_ = new_n506_ & ~new_n508_;
  assign new_n512_ = ~new_n506_ & new_n508_;
  assign new_n514_ = ~new_n510_ & ~new_n512_;
  assign new_n516_ = new_n268_ & ~new_n514_;
  assign new_n518_ = ~new_n268_ & new_n514_;
  assign new_n520_ = ~new_n516_ & ~new_n518_;
  assign new_n522_ = new_n254_ & new_n452_;
  assign new_n524_ = new_n256_ & ~new_n452_;
  assign new_n526_ = ~new_n446_ & ~new_n522_;
  assign new_n528_ = new_n524_ & ~new_n526_;
  assign new_n530_ = ~new_n524_ & new_n526_;
  assign new_n532_ = ~new_n528_ & ~new_n530_;
  assign new_n534_ = new_n268_ & ~new_n532_;
  assign new_n536_ = ~new_n268_ & new_n532_;
  assign new_n538_ = ~new_n534_ & ~new_n536_;
  assign new_n540_ = new_n256_ & new_n452_;
  assign new_n542_ = new_n258_ & ~new_n452_;
  assign new_n544_ = ~new_n446_ & ~new_n540_;
  assign new_n546_ = new_n542_ & ~new_n544_;
  assign new_n548_ = ~new_n542_ & new_n544_;
  assign new_n550_ = ~new_n546_ & ~new_n548_;
  assign new_n552_ = new_n268_ & ~new_n550_;
  assign new_n554_ = ~new_n268_ & new_n550_;
  assign new_n556_ = ~new_n552_ & ~new_n554_;
  assign new_n558_ = new_n258_ & new_n452_;
  assign new_n560_ = new_n260_ & ~new_n452_;
  assign new_n562_ = ~new_n446_ & ~new_n558_;
  assign new_n564_ = new_n560_ & ~new_n562_;
  assign new_n566_ = ~new_n560_ & new_n562_;
  assign new_n568_ = ~new_n564_ & ~new_n566_;
  assign new_n570_ = new_n268_ & ~new_n568_;
  assign new_n572_ = ~new_n268_ & new_n568_;
  assign new_n574_ = ~new_n570_ & ~new_n572_;
  assign new_n576_ = new_n260_ & new_n452_;
  assign new_n578_ = new_n262_ & ~new_n452_;
  assign new_n580_ = ~new_n446_ & ~new_n576_;
  assign new_n582_ = new_n578_ & ~new_n580_;
  assign new_n584_ = ~new_n578_ & new_n580_;
  assign new_n586_ = ~new_n582_ & ~new_n584_;
  assign new_n588_ = new_n268_ & ~new_n586_;
  assign new_n590_ = ~new_n268_ & new_n586_;
  assign new_n592_ = ~new_n588_ & ~new_n590_;
  assign new_n594_ = new_n262_ & new_n452_;
  assign new_n596_ = ~new_n446_ & ~new_n594_;
  assign new_n598_ = new_n578_ & ~new_n596_;
  assign new_n600_ = ~new_n578_ & new_n596_;
  assign new_n602_ = ~new_n598_ & ~new_n600_;
  assign new_n604_ = new_n268_ & ~new_n602_;
  assign new_n606_ = ~new_n268_ & new_n602_;
  assign new_n608_ = ~new_n604_ & ~new_n606_;
  assign new_n610_ = new_n272_ & ~new_n274_;
  assign new_n612_ = ~new_n272_ & new_n274_;
  assign new_n614_ = ~new_n610_ & ~new_n612_;
  assign new_n616_ = new_n270_ & ~new_n272_;
  assign new_n618_ = ~new_n270_ & new_n272_;
  assign new_n620_ = ~new_n616_ & ~new_n618_;
  assign new_n622_ = new_n248_ & ~new_n620_;
  assign new_n624_ = ~new_n614_ & new_n622_;
  assign new_n626_ = new_n614_ & ~new_n622_;
  assign new_n628_ = ~new_n624_ & ~new_n626_;
  assign new_n630_ = new_n272_ & ~new_n628_;
  assign new_n632_ = ~new_n272_ & new_n628_;
  assign new_n634_ = ~new_n630_ & ~new_n632_;
  assign new_n636_ = new_n248_ & new_n620_;
  assign new_n638_ = new_n250_ & ~new_n620_;
  assign new_n640_ = ~new_n614_ & ~new_n636_;
  assign new_n642_ = new_n638_ & ~new_n640_;
  assign new_n644_ = ~new_n638_ & new_n640_;
  assign new_n646_ = ~new_n642_ & ~new_n644_;
  assign new_n648_ = new_n272_ & ~new_n646_;
  assign new_n650_ = ~new_n272_ & new_n646_;
  assign new_n652_ = ~new_n648_ & ~new_n650_;
  assign new_n654_ = new_n250_ & new_n620_;
  assign new_n656_ = new_n252_ & ~new_n620_;
  assign new_n658_ = ~new_n614_ & ~new_n654_;
  assign new_n660_ = new_n656_ & ~new_n658_;
  assign new_n662_ = ~new_n656_ & new_n658_;
  assign new_n664_ = ~new_n660_ & ~new_n662_;
  assign new_n666_ = new_n272_ & ~new_n664_;
  assign new_n668_ = ~new_n272_ & new_n664_;
  assign new_n670_ = ~new_n666_ & ~new_n668_;
  assign new_n672_ = new_n252_ & new_n620_;
  assign new_n674_ = new_n254_ & ~new_n620_;
  assign new_n676_ = ~new_n614_ & ~new_n672_;
  assign new_n678_ = new_n674_ & ~new_n676_;
  assign new_n680_ = ~new_n674_ & new_n676_;
  assign new_n682_ = ~new_n678_ & ~new_n680_;
  assign new_n684_ = new_n272_ & ~new_n682_;
  assign new_n686_ = ~new_n272_ & new_n682_;
  assign new_n688_ = ~new_n684_ & ~new_n686_;
  assign new_n690_ = new_n254_ & new_n620_;
  assign new_n692_ = new_n256_ & ~new_n620_;
  assign new_n694_ = ~new_n614_ & ~new_n690_;
  assign new_n696_ = new_n692_ & ~new_n694_;
  assign new_n698_ = ~new_n692_ & new_n694_;
  assign new_n700_ = ~new_n696_ & ~new_n698_;
  assign new_n702_ = new_n272_ & ~new_n700_;
  assign new_n704_ = ~new_n272_ & new_n700_;
  assign new_n706_ = ~new_n702_ & ~new_n704_;
  assign new_n708_ = new_n256_ & new_n620_;
  assign new_n710_ = new_n258_ & ~new_n620_;
  assign new_n712_ = ~new_n614_ & ~new_n708_;
  assign new_n714_ = new_n710_ & ~new_n712_;
  assign new_n716_ = ~new_n710_ & new_n712_;
  assign new_n718_ = ~new_n714_ & ~new_n716_;
  assign new_n720_ = new_n272_ & ~new_n718_;
  assign new_n722_ = ~new_n272_ & new_n718_;
  assign new_n724_ = ~new_n720_ & ~new_n722_;
  assign new_n726_ = new_n258_ & new_n620_;
  assign new_n728_ = new_n260_ & ~new_n620_;
  assign new_n730_ = ~new_n614_ & ~new_n726_;
  assign new_n732_ = new_n728_ & ~new_n730_;
  assign new_n734_ = ~new_n728_ & new_n730_;
  assign new_n736_ = ~new_n732_ & ~new_n734_;
  assign new_n738_ = new_n272_ & ~new_n736_;
  assign new_n740_ = ~new_n272_ & new_n736_;
  assign new_n742_ = ~new_n738_ & ~new_n740_;
  assign new_n744_ = new_n260_ & new_n620_;
  assign new_n746_ = new_n262_ & ~new_n620_;
  assign new_n748_ = ~new_n614_ & ~new_n744_;
  assign new_n750_ = new_n746_ & ~new_n748_;
  assign new_n752_ = ~new_n746_ & new_n748_;
  assign new_n754_ = ~new_n750_ & ~new_n752_;
  assign new_n756_ = new_n272_ & ~new_n754_;
  assign new_n758_ = ~new_n272_ & new_n754_;
  assign new_n760_ = ~new_n756_ & ~new_n758_;
  assign new_n762_ = new_n262_ & new_n620_;
  assign new_n764_ = ~new_n614_ & ~new_n762_;
  assign new_n766_ = new_n746_ & ~new_n764_;
  assign new_n768_ = ~new_n746_ & new_n764_;
  assign new_n770_ = ~new_n766_ & ~new_n768_;
  assign new_n772_ = new_n272_ & ~new_n770_;
  assign new_n774_ = ~new_n272_ & new_n770_;
  assign new_n776_ = ~new_n772_ & ~new_n774_;
  assign new_n778_ = new_n276_ & ~new_n278_;
  assign new_n780_ = ~new_n276_ & new_n278_;
  assign new_n782_ = ~new_n778_ & ~new_n780_;
  assign new_n784_ = new_n274_ & ~new_n276_;
  assign new_n786_ = ~new_n274_ & new_n276_;
  assign new_n788_ = ~new_n784_ & ~new_n786_;
  assign new_n790_ = new_n248_ & ~new_n788_;
  assign new_n792_ = ~new_n782_ & new_n790_;
  assign new_n794_ = new_n782_ & ~new_n790_;
  assign new_n796_ = ~new_n792_ & ~new_n794_;
  assign new_n798_ = new_n276_ & ~new_n796_;
  assign new_n800_ = ~new_n276_ & new_n796_;
  assign new_n802_ = ~new_n798_ & ~new_n800_;
  assign new_n804_ = new_n248_ & new_n788_;
  assign new_n806_ = new_n250_ & ~new_n788_;
  assign new_n808_ = ~new_n782_ & ~new_n804_;
  assign new_n810_ = new_n806_ & ~new_n808_;
  assign new_n812_ = ~new_n806_ & new_n808_;
  assign new_n814_ = ~new_n810_ & ~new_n812_;
  assign new_n816_ = new_n276_ & ~new_n814_;
  assign new_n818_ = ~new_n276_ & new_n814_;
  assign new_n820_ = ~new_n816_ & ~new_n818_;
  assign new_n822_ = new_n250_ & new_n788_;
  assign new_n824_ = new_n252_ & ~new_n788_;
  assign new_n826_ = ~new_n782_ & ~new_n822_;
  assign new_n828_ = new_n824_ & ~new_n826_;
  assign new_n830_ = ~new_n824_ & new_n826_;
  assign new_n832_ = ~new_n828_ & ~new_n830_;
  assign new_n834_ = new_n276_ & ~new_n832_;
  assign new_n836_ = ~new_n276_ & new_n832_;
  assign new_n838_ = ~new_n834_ & ~new_n836_;
  assign new_n840_ = new_n252_ & new_n788_;
  assign new_n842_ = new_n254_ & ~new_n788_;
  assign new_n844_ = ~new_n782_ & ~new_n840_;
  assign new_n846_ = new_n842_ & ~new_n844_;
  assign new_n848_ = ~new_n842_ & new_n844_;
  assign new_n850_ = ~new_n846_ & ~new_n848_;
  assign new_n852_ = new_n276_ & ~new_n850_;
  assign new_n854_ = ~new_n276_ & new_n850_;
  assign new_n856_ = ~new_n852_ & ~new_n854_;
  assign new_n858_ = new_n254_ & new_n788_;
  assign new_n860_ = new_n256_ & ~new_n788_;
  assign new_n862_ = ~new_n782_ & ~new_n858_;
  assign new_n864_ = new_n860_ & ~new_n862_;
  assign new_n866_ = ~new_n860_ & new_n862_;
  assign new_n868_ = ~new_n864_ & ~new_n866_;
  assign new_n870_ = new_n276_ & ~new_n868_;
  assign new_n872_ = ~new_n276_ & new_n868_;
  assign new_n874_ = ~new_n870_ & ~new_n872_;
  assign new_n876_ = new_n256_ & new_n788_;
  assign new_n878_ = new_n258_ & ~new_n788_;
  assign new_n880_ = ~new_n782_ & ~new_n876_;
  assign new_n882_ = new_n878_ & ~new_n880_;
  assign new_n884_ = ~new_n878_ & new_n880_;
  assign new_n886_ = ~new_n882_ & ~new_n884_;
  assign new_n888_ = new_n276_ & ~new_n886_;
  assign new_n890_ = ~new_n276_ & new_n886_;
  assign new_n892_ = ~new_n888_ & ~new_n890_;
  assign new_n894_ = new_n258_ & new_n788_;
  assign new_n896_ = new_n260_ & ~new_n788_;
  assign new_n898_ = ~new_n782_ & ~new_n894_;
  assign new_n900_ = new_n896_ & ~new_n898_;
  assign new_n902_ = ~new_n896_ & new_n898_;
  assign new_n904_ = ~new_n900_ & ~new_n902_;
  assign new_n906_ = new_n276_ & ~new_n904_;
  assign new_n908_ = ~new_n276_ & new_n904_;
  assign new_n910_ = ~new_n906_ & ~new_n908_;
  assign new_n912_ = new_n260_ & new_n788_;
  assign new_n914_ = new_n262_ & ~new_n788_;
  assign new_n916_ = ~new_n782_ & ~new_n912_;
  assign new_n918_ = new_n914_ & ~new_n916_;
  assign new_n920_ = ~new_n914_ & new_n916_;
  assign new_n922_ = ~new_n918_ & ~new_n920_;
  assign new_n924_ = new_n276_ & ~new_n922_;
  assign new_n926_ = ~new_n276_ & new_n922_;
  assign new_n928_ = ~new_n924_ & ~new_n926_;
  assign new_n930_ = new_n262_ & new_n788_;
  assign new_n932_ = ~new_n782_ & ~new_n930_;
  assign new_n934_ = new_n914_ & ~new_n932_;
  assign new_n936_ = ~new_n914_ & new_n932_;
  assign new_n938_ = ~new_n934_ & ~new_n936_;
  assign new_n940_ = new_n276_ & ~new_n938_;
  assign new_n942_ = ~new_n276_ & new_n938_;
  assign new_n944_ = ~new_n940_ & ~new_n942_;
  assign \new_Multi8|y0_00_  = new_n266_;
  assign \new_Multi8|y0_01_  = new_n246_;
  assign \new_Multi8|y0_02_  = new_n270_;
  assign \new_Multi8|y0_03_  = new_n246_;
  assign \new_Multi8|y0_04_  = new_n274_;
  assign \new_Multi8|y0_05_  = new_n246_;
  assign \new_Multi8|y0_06_  = new_n278_;
  assign \new_Multi8|y0_07_  = new_n246_;
  assign \new_Multi8|y0_08_  = new_n246_;
  assign \new_Multi8|y0_09_  = new_n246_;
  assign \new_Multi8|y0_10_  = new_n246_;
  assign \new_Multi8|y0_11_  = new_n246_;
  assign \new_Multi8|y0_12_  = new_n246_;
  assign \new_Multi8|y0_13_  = new_n246_;
  assign \new_Multi8|y0_14_  = new_n246_;
  assign \new_Multi8|y0_15_  = new_n246_;
  assign \new_Multi8|y1_00_  = ~new_n298_;
  assign \new_Multi8|y1_01_  = new_n316_;
  assign \new_Multi8|y1_02_  = new_n334_;
  assign \new_Multi8|y1_03_  = new_n352_;
  assign \new_Multi8|y1_04_  = new_n370_;
  assign \new_Multi8|y1_05_  = new_n388_;
  assign \new_Multi8|y1_06_  = new_n406_;
  assign \new_Multi8|y1_07_  = new_n424_;
  assign \new_Multi8|y1_08_  = new_n440_;
  assign \new_Multi8|y1_09_  = new_n440_;
  assign \new_Multi8|y1_10_  = ~new_n440_;
  assign \new_Multi8|y1_11_  = new_n246_;
  assign \new_Multi8|y1_12_  = new_n246_;
  assign \new_Multi8|y1_13_  = new_n246_;
  assign \new_Multi8|y1_14_  = new_n246_;
  assign \new_Multi8|y1_15_  = new_n246_;
  assign \new_Multi8|y2_00_  = new_n246_;
  assign \new_Multi8|y2_01_  = new_n246_;
  assign \new_Multi8|y2_02_  = ~new_n466_;
  assign \new_Multi8|y2_03_  = new_n484_;
  assign \new_Multi8|y2_04_  = new_n502_;
  assign \new_Multi8|y2_05_  = new_n520_;
  assign \new_Multi8|y2_06_  = new_n538_;
  assign \new_Multi8|y2_07_  = new_n556_;
  assign \new_Multi8|y2_08_  = new_n574_;
  assign \new_Multi8|y2_09_  = new_n592_;
  assign \new_Multi8|y2_10_  = ~new_n608_;
  assign \new_Multi8|y2_11_  = ~new_n246_;
  assign \new_Multi8|y2_12_  = new_n246_;
  assign \new_Multi8|y2_13_  = new_n246_;
  assign \new_Multi8|y2_14_  = new_n246_;
  assign \new_Multi8|y2_15_  = new_n246_;
  assign \new_Multi8|y3_00_  = new_n246_;
  assign \new_Multi8|y3_01_  = new_n246_;
  assign \new_Multi8|y3_02_  = new_n246_;
  assign \new_Multi8|y3_03_  = new_n246_;
  assign \new_Multi8|y3_04_  = ~new_n634_;
  assign \new_Multi8|y3_05_  = new_n652_;
  assign \new_Multi8|y3_06_  = new_n670_;
  assign \new_Multi8|y3_07_  = new_n688_;
  assign \new_Multi8|y3_08_  = new_n706_;
  assign \new_Multi8|y3_09_  = new_n724_;
  assign \new_Multi8|y3_10_  = new_n742_;
  assign \new_Multi8|y3_11_  = new_n760_;
  assign \new_Multi8|y3_12_  = ~new_n776_;
  assign \new_Multi8|y3_13_  = ~new_n246_;
  assign \new_Multi8|y3_14_  = new_n246_;
  assign \new_Multi8|y3_15_  = new_n246_;
  assign \new_Multi8|y4_00_  = new_n246_;
  assign \new_Multi8|y4_01_  = new_n246_;
  assign \new_Multi8|y4_02_  = new_n246_;
  assign \new_Multi8|y4_03_  = new_n246_;
  assign \new_Multi8|y4_04_  = new_n246_;
  assign \new_Multi8|y4_05_  = new_n246_;
  assign \new_Multi8|y4_06_  = ~new_n802_;
  assign \new_Multi8|y4_07_  = new_n820_;
  assign \new_Multi8|y4_08_  = new_n838_;
  assign \new_Multi8|y4_09_  = new_n856_;
  assign \new_Multi8|y4_10_  = new_n874_;
  assign \new_Multi8|y4_11_  = new_n892_;
  assign \new_Multi8|y4_12_  = new_n910_;
  assign \new_Multi8|y4_13_  = new_n928_;
  assign \new_Multi8|y4_14_  = ~new_n944_;
  assign \new_Multi8|y4_15_  = ~new_n246_;
  assign \new_Multi8|x0_00_  = 1'b0;
  assign \new_Multi8|x0_01_  = 1'b0;
  assign \new_Multi8|x0_02_  = 1'b0;
  assign \new_Multi8|x0_03_  = 1'b0;
  assign \new_Multi8|x0_04_  = 1'b0;
  assign \new_Multi8|x0_05_  = 1'b0;
  assign \new_Multi8|x0_06_  = 1'b0;
  assign \new_Multi8|x0_07_  = 1'b0;
  assign \new_Multi8|x0_08_  = 1'b0;
  assign \new_Multi8|x0_09_  = 1'b0;
  assign \new_Multi8|x0_10_  = 1'b0;
  assign \new_Multi8|x0_11_  = 1'b0;
  assign \new_Multi8|x0_12_  = 1'b0;
  assign \new_Multi8|x0_13_  = 1'b0;
  assign \new_Multi8|x0_14_  = 1'b0;
  assign \new_Multi8|x0_15_  = 1'b0;
  assign m00 = \new_Multi8|x5_00_ ;
  assign m01 = \new_Multi8|x5_01_ ;
  assign m02 = \new_Multi8|x5_02_ ;
  assign m03 = \new_Multi8|x5_03_ ;
  assign m04 = \new_Multi8|x5_04_ ;
  assign m05 = \new_Multi8|x5_05_ ;
  assign m06 = \new_Multi8|x5_06_ ;
  assign m07 = \new_Multi8|x5_07_ ;
  assign m08 = \new_Multi8|x5_08_ ;
  assign m09 = \new_Multi8|x5_09_ ;
  assign m10 = \new_Multi8|x5_10_ ;
  assign m11 = \new_Multi8|x5_11_ ;
  assign m12 = \new_Multi8|x5_12_ ;
  assign m13 = \new_Multi8|x5_13_ ;
  assign m14 = \new_Multi8|x5_14_ ;
  assign m15 = \new_Multi8|x5_15_ ;
  assign \new_Multi8|ADD16(1)|c_  = 1'b0;
  assign new_n1075_ = \new_Multi8|x0_00_  & \new_Multi8|y0_00_ ;
  assign new_n1077_ = ~\new_Multi8|x0_00_  & ~\new_Multi8|y0_00_ ;
  assign new_n1079_ = ~new_n1075_ & ~new_n1077_;
  assign new_n1081_ = \new_Multi8|ADD16(1)|c_  & new_n1079_;
  assign new_n1083_ = ~\new_Multi8|ADD16(1)|c_  & ~new_n1079_;
  assign \new_Multi8|x1_00_  = ~new_n1081_ & ~new_n1083_;
  assign \new_Multi8|ADD16(1)|00_  = new_n1075_ | new_n1081_;
  assign new_n1087_ = \new_Multi8|x0_01_  & \new_Multi8|y0_01_ ;
  assign new_n1089_ = ~\new_Multi8|x0_01_  & ~\new_Multi8|y0_01_ ;
  assign new_n1091_ = ~new_n1087_ & ~new_n1089_;
  assign new_n1093_ = \new_Multi8|ADD16(1)|00_  & new_n1091_;
  assign new_n1095_ = ~\new_Multi8|ADD16(1)|00_  & ~new_n1091_;
  assign \new_Multi8|x1_01_  = ~new_n1093_ & ~new_n1095_;
  assign \new_Multi8|ADD16(1)|01_  = new_n1087_ | new_n1093_;
  assign new_n1099_ = \new_Multi8|x0_02_  & \new_Multi8|y0_02_ ;
  assign new_n1101_ = ~\new_Multi8|x0_02_  & ~\new_Multi8|y0_02_ ;
  assign new_n1103_ = ~new_n1099_ & ~new_n1101_;
  assign new_n1105_ = \new_Multi8|ADD16(1)|01_  & new_n1103_;
  assign new_n1107_ = ~\new_Multi8|ADD16(1)|01_  & ~new_n1103_;
  assign \new_Multi8|x1_02_  = ~new_n1105_ & ~new_n1107_;
  assign \new_Multi8|ADD16(1)|02_  = new_n1099_ | new_n1105_;
  assign new_n1111_ = \new_Multi8|x0_03_  & \new_Multi8|y0_03_ ;
  assign new_n1113_ = ~\new_Multi8|x0_03_  & ~\new_Multi8|y0_03_ ;
  assign new_n1115_ = ~new_n1111_ & ~new_n1113_;
  assign new_n1117_ = \new_Multi8|ADD16(1)|02_  & new_n1115_;
  assign new_n1119_ = ~\new_Multi8|ADD16(1)|02_  & ~new_n1115_;
  assign \new_Multi8|x1_03_  = ~new_n1117_ & ~new_n1119_;
  assign \new_Multi8|ADD16(1)|03_  = new_n1111_ | new_n1117_;
  assign new_n1123_ = \new_Multi8|x0_04_  & \new_Multi8|y0_04_ ;
  assign new_n1125_ = ~\new_Multi8|x0_04_  & ~\new_Multi8|y0_04_ ;
  assign new_n1127_ = ~new_n1123_ & ~new_n1125_;
  assign new_n1129_ = \new_Multi8|ADD16(1)|03_  & new_n1127_;
  assign new_n1131_ = ~\new_Multi8|ADD16(1)|03_  & ~new_n1127_;
  assign \new_Multi8|x1_04_  = ~new_n1129_ & ~new_n1131_;
  assign \new_Multi8|ADD16(1)|04_  = new_n1123_ | new_n1129_;
  assign new_n1135_ = \new_Multi8|x0_05_  & \new_Multi8|y0_05_ ;
  assign new_n1137_ = ~\new_Multi8|x0_05_  & ~\new_Multi8|y0_05_ ;
  assign new_n1139_ = ~new_n1135_ & ~new_n1137_;
  assign new_n1141_ = \new_Multi8|ADD16(1)|04_  & new_n1139_;
  assign new_n1143_ = ~\new_Multi8|ADD16(1)|04_  & ~new_n1139_;
  assign \new_Multi8|x1_05_  = ~new_n1141_ & ~new_n1143_;
  assign \new_Multi8|ADD16(1)|05_  = new_n1135_ | new_n1141_;
  assign new_n1147_ = \new_Multi8|x0_06_  & \new_Multi8|y0_06_ ;
  assign new_n1149_ = ~\new_Multi8|x0_06_  & ~\new_Multi8|y0_06_ ;
  assign new_n1151_ = ~new_n1147_ & ~new_n1149_;
  assign new_n1153_ = \new_Multi8|ADD16(1)|05_  & new_n1151_;
  assign new_n1155_ = ~\new_Multi8|ADD16(1)|05_  & ~new_n1151_;
  assign \new_Multi8|x1_06_  = ~new_n1153_ & ~new_n1155_;
  assign \new_Multi8|ADD16(1)|06_  = new_n1147_ | new_n1153_;
  assign new_n1159_ = \new_Multi8|x0_07_  & \new_Multi8|y0_07_ ;
  assign new_n1161_ = ~\new_Multi8|x0_07_  & ~\new_Multi8|y0_07_ ;
  assign new_n1163_ = ~new_n1159_ & ~new_n1161_;
  assign new_n1165_ = \new_Multi8|ADD16(1)|06_  & new_n1163_;
  assign new_n1167_ = ~\new_Multi8|ADD16(1)|06_  & ~new_n1163_;
  assign \new_Multi8|x1_07_  = ~new_n1165_ & ~new_n1167_;
  assign \new_Multi8|ADD16(1)|07_  = new_n1159_ | new_n1165_;
  assign new_n1171_ = \new_Multi8|x0_08_  & \new_Multi8|y0_08_ ;
  assign new_n1173_ = ~\new_Multi8|x0_08_  & ~\new_Multi8|y0_08_ ;
  assign new_n1175_ = ~new_n1171_ & ~new_n1173_;
  assign new_n1177_ = \new_Multi8|ADD16(1)|07_  & new_n1175_;
  assign new_n1179_ = ~\new_Multi8|ADD16(1)|07_  & ~new_n1175_;
  assign \new_Multi8|x1_08_  = ~new_n1177_ & ~new_n1179_;
  assign \new_Multi8|ADD16(1)|08_  = new_n1171_ | new_n1177_;
  assign new_n1183_ = \new_Multi8|x0_09_  & \new_Multi8|y0_09_ ;
  assign new_n1185_ = ~\new_Multi8|x0_09_  & ~\new_Multi8|y0_09_ ;
  assign new_n1187_ = ~new_n1183_ & ~new_n1185_;
  assign new_n1189_ = \new_Multi8|ADD16(1)|08_  & new_n1187_;
  assign new_n1191_ = ~\new_Multi8|ADD16(1)|08_  & ~new_n1187_;
  assign \new_Multi8|x1_09_  = ~new_n1189_ & ~new_n1191_;
  assign \new_Multi8|ADD16(1)|09_  = new_n1183_ | new_n1189_;
  assign new_n1195_ = \new_Multi8|x0_10_  & \new_Multi8|y0_10_ ;
  assign new_n1197_ = ~\new_Multi8|x0_10_  & ~\new_Multi8|y0_10_ ;
  assign new_n1199_ = ~new_n1195_ & ~new_n1197_;
  assign new_n1201_ = \new_Multi8|ADD16(1)|09_  & new_n1199_;
  assign new_n1203_ = ~\new_Multi8|ADD16(1)|09_  & ~new_n1199_;
  assign \new_Multi8|x1_10_  = ~new_n1201_ & ~new_n1203_;
  assign \new_Multi8|ADD16(1)|10_  = new_n1195_ | new_n1201_;
  assign new_n1207_ = \new_Multi8|x0_11_  & \new_Multi8|y0_11_ ;
  assign new_n1209_ = ~\new_Multi8|x0_11_  & ~\new_Multi8|y0_11_ ;
  assign new_n1211_ = ~new_n1207_ & ~new_n1209_;
  assign new_n1213_ = \new_Multi8|ADD16(1)|10_  & new_n1211_;
  assign new_n1215_ = ~\new_Multi8|ADD16(1)|10_  & ~new_n1211_;
  assign \new_Multi8|x1_11_  = ~new_n1213_ & ~new_n1215_;
  assign \new_Multi8|ADD16(1)|11_  = new_n1207_ | new_n1213_;
  assign new_n1219_ = \new_Multi8|x0_12_  & \new_Multi8|y0_12_ ;
  assign new_n1221_ = ~\new_Multi8|x0_12_  & ~\new_Multi8|y0_12_ ;
  assign new_n1223_ = ~new_n1219_ & ~new_n1221_;
  assign new_n1225_ = \new_Multi8|ADD16(1)|11_  & new_n1223_;
  assign new_n1227_ = ~\new_Multi8|ADD16(1)|11_  & ~new_n1223_;
  assign \new_Multi8|x1_12_  = ~new_n1225_ & ~new_n1227_;
  assign \new_Multi8|ADD16(1)|12_  = new_n1219_ | new_n1225_;
  assign new_n1231_ = \new_Multi8|x0_13_  & \new_Multi8|y0_13_ ;
  assign new_n1233_ = ~\new_Multi8|x0_13_  & ~\new_Multi8|y0_13_ ;
  assign new_n1235_ = ~new_n1231_ & ~new_n1233_;
  assign new_n1237_ = \new_Multi8|ADD16(1)|12_  & new_n1235_;
  assign new_n1239_ = ~\new_Multi8|ADD16(1)|12_  & ~new_n1235_;
  assign \new_Multi8|x1_13_  = ~new_n1237_ & ~new_n1239_;
  assign \new_Multi8|ADD16(1)|13_  = new_n1231_ | new_n1237_;
  assign new_n1243_ = \new_Multi8|x0_14_  & \new_Multi8|y0_14_ ;
  assign new_n1245_ = ~\new_Multi8|x0_14_  & ~\new_Multi8|y0_14_ ;
  assign new_n1247_ = ~new_n1243_ & ~new_n1245_;
  assign new_n1249_ = \new_Multi8|ADD16(1)|13_  & new_n1247_;
  assign new_n1251_ = ~\new_Multi8|ADD16(1)|13_  & ~new_n1247_;
  assign \new_Multi8|x1_14_  = ~new_n1249_ & ~new_n1251_;
  assign \new_Multi8|ADD16(1)|14_  = new_n1243_ | new_n1249_;
  assign new_n1255_ = \new_Multi8|x0_15_  & \new_Multi8|y0_15_ ;
  assign new_n1257_ = ~\new_Multi8|x0_15_  & ~\new_Multi8|y0_15_ ;
  assign new_n1259_ = ~new_n1255_ & ~new_n1257_;
  assign new_n1261_ = \new_Multi8|ADD16(1)|14_  & new_n1259_;
  assign new_n1263_ = ~\new_Multi8|ADD16(1)|14_  & ~new_n1259_;
  assign \new_Multi8|x1_15_  = ~new_n1261_ & ~new_n1263_;
  assign \new_Multi8|ADD16(18)|c_  = 1'b0;
  assign new_n1284_ = \new_Multi8|x1_00_  & \new_Multi8|y1_00_ ;
  assign new_n1286_ = ~\new_Multi8|x1_00_  & ~\new_Multi8|y1_00_ ;
  assign new_n1288_ = ~new_n1284_ & ~new_n1286_;
  assign new_n1290_ = \new_Multi8|ADD16(18)|c_  & new_n1288_;
  assign new_n1292_ = ~\new_Multi8|ADD16(18)|c_  & ~new_n1288_;
  assign \new_Multi8|x2_00_  = ~new_n1290_ & ~new_n1292_;
  assign \new_Multi8|ADD16(18)|00_  = new_n1284_ | new_n1290_;
  assign new_n1296_ = \new_Multi8|x1_01_  & \new_Multi8|y1_01_ ;
  assign new_n1298_ = ~\new_Multi8|x1_01_  & ~\new_Multi8|y1_01_ ;
  assign new_n1300_ = ~new_n1296_ & ~new_n1298_;
  assign new_n1302_ = \new_Multi8|ADD16(18)|00_  & new_n1300_;
  assign new_n1304_ = ~\new_Multi8|ADD16(18)|00_  & ~new_n1300_;
  assign \new_Multi8|x2_01_  = ~new_n1302_ & ~new_n1304_;
  assign \new_Multi8|ADD16(18)|01_  = new_n1296_ | new_n1302_;
  assign new_n1308_ = \new_Multi8|x1_02_  & \new_Multi8|y1_02_ ;
  assign new_n1310_ = ~\new_Multi8|x1_02_  & ~\new_Multi8|y1_02_ ;
  assign new_n1312_ = ~new_n1308_ & ~new_n1310_;
  assign new_n1314_ = \new_Multi8|ADD16(18)|01_  & new_n1312_;
  assign new_n1316_ = ~\new_Multi8|ADD16(18)|01_  & ~new_n1312_;
  assign \new_Multi8|x2_02_  = ~new_n1314_ & ~new_n1316_;
  assign \new_Multi8|ADD16(18)|02_  = new_n1308_ | new_n1314_;
  assign new_n1320_ = \new_Multi8|x1_03_  & \new_Multi8|y1_03_ ;
  assign new_n1322_ = ~\new_Multi8|x1_03_  & ~\new_Multi8|y1_03_ ;
  assign new_n1324_ = ~new_n1320_ & ~new_n1322_;
  assign new_n1326_ = \new_Multi8|ADD16(18)|02_  & new_n1324_;
  assign new_n1328_ = ~\new_Multi8|ADD16(18)|02_  & ~new_n1324_;
  assign \new_Multi8|x2_03_  = ~new_n1326_ & ~new_n1328_;
  assign \new_Multi8|ADD16(18)|03_  = new_n1320_ | new_n1326_;
  assign new_n1332_ = \new_Multi8|x1_04_  & \new_Multi8|y1_04_ ;
  assign new_n1334_ = ~\new_Multi8|x1_04_  & ~\new_Multi8|y1_04_ ;
  assign new_n1336_ = ~new_n1332_ & ~new_n1334_;
  assign new_n1338_ = \new_Multi8|ADD16(18)|03_  & new_n1336_;
  assign new_n1340_ = ~\new_Multi8|ADD16(18)|03_  & ~new_n1336_;
  assign \new_Multi8|x2_04_  = ~new_n1338_ & ~new_n1340_;
  assign \new_Multi8|ADD16(18)|04_  = new_n1332_ | new_n1338_;
  assign new_n1344_ = \new_Multi8|x1_05_  & \new_Multi8|y1_05_ ;
  assign new_n1346_ = ~\new_Multi8|x1_05_  & ~\new_Multi8|y1_05_ ;
  assign new_n1348_ = ~new_n1344_ & ~new_n1346_;
  assign new_n1350_ = \new_Multi8|ADD16(18)|04_  & new_n1348_;
  assign new_n1352_ = ~\new_Multi8|ADD16(18)|04_  & ~new_n1348_;
  assign \new_Multi8|x2_05_  = ~new_n1350_ & ~new_n1352_;
  assign \new_Multi8|ADD16(18)|05_  = new_n1344_ | new_n1350_;
  assign new_n1356_ = \new_Multi8|x1_06_  & \new_Multi8|y1_06_ ;
  assign new_n1358_ = ~\new_Multi8|x1_06_  & ~\new_Multi8|y1_06_ ;
  assign new_n1360_ = ~new_n1356_ & ~new_n1358_;
  assign new_n1362_ = \new_Multi8|ADD16(18)|05_  & new_n1360_;
  assign new_n1364_ = ~\new_Multi8|ADD16(18)|05_  & ~new_n1360_;
  assign \new_Multi8|x2_06_  = ~new_n1362_ & ~new_n1364_;
  assign \new_Multi8|ADD16(18)|06_  = new_n1356_ | new_n1362_;
  assign new_n1368_ = \new_Multi8|x1_07_  & \new_Multi8|y1_07_ ;
  assign new_n1370_ = ~\new_Multi8|x1_07_  & ~\new_Multi8|y1_07_ ;
  assign new_n1372_ = ~new_n1368_ & ~new_n1370_;
  assign new_n1374_ = \new_Multi8|ADD16(18)|06_  & new_n1372_;
  assign new_n1376_ = ~\new_Multi8|ADD16(18)|06_  & ~new_n1372_;
  assign \new_Multi8|x2_07_  = ~new_n1374_ & ~new_n1376_;
  assign \new_Multi8|ADD16(18)|07_  = new_n1368_ | new_n1374_;
  assign new_n1380_ = \new_Multi8|x1_08_  & \new_Multi8|y1_08_ ;
  assign new_n1382_ = ~\new_Multi8|x1_08_  & ~\new_Multi8|y1_08_ ;
  assign new_n1384_ = ~new_n1380_ & ~new_n1382_;
  assign new_n1386_ = \new_Multi8|ADD16(18)|07_  & new_n1384_;
  assign new_n1388_ = ~\new_Multi8|ADD16(18)|07_  & ~new_n1384_;
  assign \new_Multi8|x2_08_  = ~new_n1386_ & ~new_n1388_;
  assign \new_Multi8|ADD16(18)|08_  = new_n1380_ | new_n1386_;
  assign new_n1392_ = \new_Multi8|x1_09_  & \new_Multi8|y1_09_ ;
  assign new_n1394_ = ~\new_Multi8|x1_09_  & ~\new_Multi8|y1_09_ ;
  assign new_n1396_ = ~new_n1392_ & ~new_n1394_;
  assign new_n1398_ = \new_Multi8|ADD16(18)|08_  & new_n1396_;
  assign new_n1400_ = ~\new_Multi8|ADD16(18)|08_  & ~new_n1396_;
  assign \new_Multi8|x2_09_  = ~new_n1398_ & ~new_n1400_;
  assign \new_Multi8|ADD16(18)|09_  = new_n1392_ | new_n1398_;
  assign new_n1404_ = \new_Multi8|x1_10_  & \new_Multi8|y1_10_ ;
  assign new_n1406_ = ~\new_Multi8|x1_10_  & ~\new_Multi8|y1_10_ ;
  assign new_n1408_ = ~new_n1404_ & ~new_n1406_;
  assign new_n1410_ = \new_Multi8|ADD16(18)|09_  & new_n1408_;
  assign new_n1412_ = ~\new_Multi8|ADD16(18)|09_  & ~new_n1408_;
  assign \new_Multi8|x2_10_  = ~new_n1410_ & ~new_n1412_;
  assign \new_Multi8|ADD16(18)|10_  = new_n1404_ | new_n1410_;
  assign new_n1416_ = \new_Multi8|x1_11_  & \new_Multi8|y1_11_ ;
  assign new_n1418_ = ~\new_Multi8|x1_11_  & ~\new_Multi8|y1_11_ ;
  assign new_n1420_ = ~new_n1416_ & ~new_n1418_;
  assign new_n1422_ = \new_Multi8|ADD16(18)|10_  & new_n1420_;
  assign new_n1424_ = ~\new_Multi8|ADD16(18)|10_  & ~new_n1420_;
  assign \new_Multi8|x2_11_  = ~new_n1422_ & ~new_n1424_;
  assign \new_Multi8|ADD16(18)|11_  = new_n1416_ | new_n1422_;
  assign new_n1428_ = \new_Multi8|x1_12_  & \new_Multi8|y1_12_ ;
  assign new_n1430_ = ~\new_Multi8|x1_12_  & ~\new_Multi8|y1_12_ ;
  assign new_n1432_ = ~new_n1428_ & ~new_n1430_;
  assign new_n1434_ = \new_Multi8|ADD16(18)|11_  & new_n1432_;
  assign new_n1436_ = ~\new_Multi8|ADD16(18)|11_  & ~new_n1432_;
  assign \new_Multi8|x2_12_  = ~new_n1434_ & ~new_n1436_;
  assign \new_Multi8|ADD16(18)|12_  = new_n1428_ | new_n1434_;
  assign new_n1440_ = \new_Multi8|x1_13_  & \new_Multi8|y1_13_ ;
  assign new_n1442_ = ~\new_Multi8|x1_13_  & ~\new_Multi8|y1_13_ ;
  assign new_n1444_ = ~new_n1440_ & ~new_n1442_;
  assign new_n1446_ = \new_Multi8|ADD16(18)|12_  & new_n1444_;
  assign new_n1448_ = ~\new_Multi8|ADD16(18)|12_  & ~new_n1444_;
  assign \new_Multi8|x2_13_  = ~new_n1446_ & ~new_n1448_;
  assign \new_Multi8|ADD16(18)|13_  = new_n1440_ | new_n1446_;
  assign new_n1452_ = \new_Multi8|x1_14_  & \new_Multi8|y1_14_ ;
  assign new_n1454_ = ~\new_Multi8|x1_14_  & ~\new_Multi8|y1_14_ ;
  assign new_n1456_ = ~new_n1452_ & ~new_n1454_;
  assign new_n1458_ = \new_Multi8|ADD16(18)|13_  & new_n1456_;
  assign new_n1460_ = ~\new_Multi8|ADD16(18)|13_  & ~new_n1456_;
  assign \new_Multi8|x2_14_  = ~new_n1458_ & ~new_n1460_;
  assign \new_Multi8|ADD16(18)|14_  = new_n1452_ | new_n1458_;
  assign new_n1464_ = \new_Multi8|x1_15_  & \new_Multi8|y1_15_ ;
  assign new_n1466_ = ~\new_Multi8|x1_15_  & ~\new_Multi8|y1_15_ ;
  assign new_n1468_ = ~new_n1464_ & ~new_n1466_;
  assign new_n1470_ = \new_Multi8|ADD16(18)|14_  & new_n1468_;
  assign new_n1472_ = ~\new_Multi8|ADD16(18)|14_  & ~new_n1468_;
  assign \new_Multi8|x2_15_  = ~new_n1470_ & ~new_n1472_;
  assign \new_Multi8|ADD16(35)|c_  = 1'b0;
  assign new_n1493_ = \new_Multi8|x2_00_  & \new_Multi8|y2_00_ ;
  assign new_n1495_ = ~\new_Multi8|x2_00_  & ~\new_Multi8|y2_00_ ;
  assign new_n1497_ = ~new_n1493_ & ~new_n1495_;
  assign new_n1499_ = \new_Multi8|ADD16(35)|c_  & new_n1497_;
  assign new_n1501_ = ~\new_Multi8|ADD16(35)|c_  & ~new_n1497_;
  assign \new_Multi8|x3_00_  = ~new_n1499_ & ~new_n1501_;
  assign \new_Multi8|ADD16(35)|00_  = new_n1493_ | new_n1499_;
  assign new_n1505_ = \new_Multi8|x2_01_  & \new_Multi8|y2_01_ ;
  assign new_n1507_ = ~\new_Multi8|x2_01_  & ~\new_Multi8|y2_01_ ;
  assign new_n1509_ = ~new_n1505_ & ~new_n1507_;
  assign new_n1511_ = \new_Multi8|ADD16(35)|00_  & new_n1509_;
  assign new_n1513_ = ~\new_Multi8|ADD16(35)|00_  & ~new_n1509_;
  assign \new_Multi8|x3_01_  = ~new_n1511_ & ~new_n1513_;
  assign \new_Multi8|ADD16(35)|01_  = new_n1505_ | new_n1511_;
  assign new_n1517_ = \new_Multi8|x2_02_  & \new_Multi8|y2_02_ ;
  assign new_n1519_ = ~\new_Multi8|x2_02_  & ~\new_Multi8|y2_02_ ;
  assign new_n1521_ = ~new_n1517_ & ~new_n1519_;
  assign new_n1523_ = \new_Multi8|ADD16(35)|01_  & new_n1521_;
  assign new_n1525_ = ~\new_Multi8|ADD16(35)|01_  & ~new_n1521_;
  assign \new_Multi8|x3_02_  = ~new_n1523_ & ~new_n1525_;
  assign \new_Multi8|ADD16(35)|02_  = new_n1517_ | new_n1523_;
  assign new_n1529_ = \new_Multi8|x2_03_  & \new_Multi8|y2_03_ ;
  assign new_n1531_ = ~\new_Multi8|x2_03_  & ~\new_Multi8|y2_03_ ;
  assign new_n1533_ = ~new_n1529_ & ~new_n1531_;
  assign new_n1535_ = \new_Multi8|ADD16(35)|02_  & new_n1533_;
  assign new_n1537_ = ~\new_Multi8|ADD16(35)|02_  & ~new_n1533_;
  assign \new_Multi8|x3_03_  = ~new_n1535_ & ~new_n1537_;
  assign \new_Multi8|ADD16(35)|03_  = new_n1529_ | new_n1535_;
  assign new_n1541_ = \new_Multi8|x2_04_  & \new_Multi8|y2_04_ ;
  assign new_n1543_ = ~\new_Multi8|x2_04_  & ~\new_Multi8|y2_04_ ;
  assign new_n1545_ = ~new_n1541_ & ~new_n1543_;
  assign new_n1547_ = \new_Multi8|ADD16(35)|03_  & new_n1545_;
  assign new_n1549_ = ~\new_Multi8|ADD16(35)|03_  & ~new_n1545_;
  assign \new_Multi8|x3_04_  = ~new_n1547_ & ~new_n1549_;
  assign \new_Multi8|ADD16(35)|04_  = new_n1541_ | new_n1547_;
  assign new_n1553_ = \new_Multi8|x2_05_  & \new_Multi8|y2_05_ ;
  assign new_n1555_ = ~\new_Multi8|x2_05_  & ~\new_Multi8|y2_05_ ;
  assign new_n1557_ = ~new_n1553_ & ~new_n1555_;
  assign new_n1559_ = \new_Multi8|ADD16(35)|04_  & new_n1557_;
  assign new_n1561_ = ~\new_Multi8|ADD16(35)|04_  & ~new_n1557_;
  assign \new_Multi8|x3_05_  = ~new_n1559_ & ~new_n1561_;
  assign \new_Multi8|ADD16(35)|05_  = new_n1553_ | new_n1559_;
  assign new_n1565_ = \new_Multi8|x2_06_  & \new_Multi8|y2_06_ ;
  assign new_n1567_ = ~\new_Multi8|x2_06_  & ~\new_Multi8|y2_06_ ;
  assign new_n1569_ = ~new_n1565_ & ~new_n1567_;
  assign new_n1571_ = \new_Multi8|ADD16(35)|05_  & new_n1569_;
  assign new_n1573_ = ~\new_Multi8|ADD16(35)|05_  & ~new_n1569_;
  assign \new_Multi8|x3_06_  = ~new_n1571_ & ~new_n1573_;
  assign \new_Multi8|ADD16(35)|06_  = new_n1565_ | new_n1571_;
  assign new_n1577_ = \new_Multi8|x2_07_  & \new_Multi8|y2_07_ ;
  assign new_n1579_ = ~\new_Multi8|x2_07_  & ~\new_Multi8|y2_07_ ;
  assign new_n1581_ = ~new_n1577_ & ~new_n1579_;
  assign new_n1583_ = \new_Multi8|ADD16(35)|06_  & new_n1581_;
  assign new_n1585_ = ~\new_Multi8|ADD16(35)|06_  & ~new_n1581_;
  assign \new_Multi8|x3_07_  = ~new_n1583_ & ~new_n1585_;
  assign \new_Multi8|ADD16(35)|07_  = new_n1577_ | new_n1583_;
  assign new_n1589_ = \new_Multi8|x2_08_  & \new_Multi8|y2_08_ ;
  assign new_n1591_ = ~\new_Multi8|x2_08_  & ~\new_Multi8|y2_08_ ;
  assign new_n1593_ = ~new_n1589_ & ~new_n1591_;
  assign new_n1595_ = \new_Multi8|ADD16(35)|07_  & new_n1593_;
  assign new_n1597_ = ~\new_Multi8|ADD16(35)|07_  & ~new_n1593_;
  assign \new_Multi8|x3_08_  = ~new_n1595_ & ~new_n1597_;
  assign \new_Multi8|ADD16(35)|08_  = new_n1589_ | new_n1595_;
  assign new_n1601_ = \new_Multi8|x2_09_  & \new_Multi8|y2_09_ ;
  assign new_n1603_ = ~\new_Multi8|x2_09_  & ~\new_Multi8|y2_09_ ;
  assign new_n1605_ = ~new_n1601_ & ~new_n1603_;
  assign new_n1607_ = \new_Multi8|ADD16(35)|08_  & new_n1605_;
  assign new_n1609_ = ~\new_Multi8|ADD16(35)|08_  & ~new_n1605_;
  assign \new_Multi8|x3_09_  = ~new_n1607_ & ~new_n1609_;
  assign \new_Multi8|ADD16(35)|09_  = new_n1601_ | new_n1607_;
  assign new_n1613_ = \new_Multi8|x2_10_  & \new_Multi8|y2_10_ ;
  assign new_n1615_ = ~\new_Multi8|x2_10_  & ~\new_Multi8|y2_10_ ;
  assign new_n1617_ = ~new_n1613_ & ~new_n1615_;
  assign new_n1619_ = \new_Multi8|ADD16(35)|09_  & new_n1617_;
  assign new_n1621_ = ~\new_Multi8|ADD16(35)|09_  & ~new_n1617_;
  assign \new_Multi8|x3_10_  = ~new_n1619_ & ~new_n1621_;
  assign \new_Multi8|ADD16(35)|10_  = new_n1613_ | new_n1619_;
  assign new_n1625_ = \new_Multi8|x2_11_  & \new_Multi8|y2_11_ ;
  assign new_n1627_ = ~\new_Multi8|x2_11_  & ~\new_Multi8|y2_11_ ;
  assign new_n1629_ = ~new_n1625_ & ~new_n1627_;
  assign new_n1631_ = \new_Multi8|ADD16(35)|10_  & new_n1629_;
  assign new_n1633_ = ~\new_Multi8|ADD16(35)|10_  & ~new_n1629_;
  assign \new_Multi8|x3_11_  = ~new_n1631_ & ~new_n1633_;
  assign \new_Multi8|ADD16(35)|11_  = new_n1625_ | new_n1631_;
  assign new_n1637_ = \new_Multi8|x2_12_  & \new_Multi8|y2_12_ ;
  assign new_n1639_ = ~\new_Multi8|x2_12_  & ~\new_Multi8|y2_12_ ;
  assign new_n1641_ = ~new_n1637_ & ~new_n1639_;
  assign new_n1643_ = \new_Multi8|ADD16(35)|11_  & new_n1641_;
  assign new_n1645_ = ~\new_Multi8|ADD16(35)|11_  & ~new_n1641_;
  assign \new_Multi8|x3_12_  = ~new_n1643_ & ~new_n1645_;
  assign \new_Multi8|ADD16(35)|12_  = new_n1637_ | new_n1643_;
  assign new_n1649_ = \new_Multi8|x2_13_  & \new_Multi8|y2_13_ ;
  assign new_n1651_ = ~\new_Multi8|x2_13_  & ~\new_Multi8|y2_13_ ;
  assign new_n1653_ = ~new_n1649_ & ~new_n1651_;
  assign new_n1655_ = \new_Multi8|ADD16(35)|12_  & new_n1653_;
  assign new_n1657_ = ~\new_Multi8|ADD16(35)|12_  & ~new_n1653_;
  assign \new_Multi8|x3_13_  = ~new_n1655_ & ~new_n1657_;
  assign \new_Multi8|ADD16(35)|13_  = new_n1649_ | new_n1655_;
  assign new_n1661_ = \new_Multi8|x2_14_  & \new_Multi8|y2_14_ ;
  assign new_n1663_ = ~\new_Multi8|x2_14_  & ~\new_Multi8|y2_14_ ;
  assign new_n1665_ = ~new_n1661_ & ~new_n1663_;
  assign new_n1667_ = \new_Multi8|ADD16(35)|13_  & new_n1665_;
  assign new_n1669_ = ~\new_Multi8|ADD16(35)|13_  & ~new_n1665_;
  assign \new_Multi8|x3_14_  = ~new_n1667_ & ~new_n1669_;
  assign \new_Multi8|ADD16(35)|14_  = new_n1661_ | new_n1667_;
  assign new_n1673_ = \new_Multi8|x2_15_  & \new_Multi8|y2_15_ ;
  assign new_n1675_ = ~\new_Multi8|x2_15_  & ~\new_Multi8|y2_15_ ;
  assign new_n1677_ = ~new_n1673_ & ~new_n1675_;
  assign new_n1679_ = \new_Multi8|ADD16(35)|14_  & new_n1677_;
  assign new_n1681_ = ~\new_Multi8|ADD16(35)|14_  & ~new_n1677_;
  assign \new_Multi8|x3_15_  = ~new_n1679_ & ~new_n1681_;
  assign \new_Multi8|ADD16(52)|c_  = 1'b0;
  assign new_n1702_ = \new_Multi8|x3_00_  & \new_Multi8|y3_00_ ;
  assign new_n1704_ = ~\new_Multi8|x3_00_  & ~\new_Multi8|y3_00_ ;
  assign new_n1706_ = ~new_n1702_ & ~new_n1704_;
  assign new_n1708_ = \new_Multi8|ADD16(52)|c_  & new_n1706_;
  assign new_n1710_ = ~\new_Multi8|ADD16(52)|c_  & ~new_n1706_;
  assign \new_Multi8|x4_00_  = ~new_n1708_ & ~new_n1710_;
  assign \new_Multi8|ADD16(52)|00_  = new_n1702_ | new_n1708_;
  assign new_n1714_ = \new_Multi8|x3_01_  & \new_Multi8|y3_01_ ;
  assign new_n1716_ = ~\new_Multi8|x3_01_  & ~\new_Multi8|y3_01_ ;
  assign new_n1718_ = ~new_n1714_ & ~new_n1716_;
  assign new_n1720_ = \new_Multi8|ADD16(52)|00_  & new_n1718_;
  assign new_n1722_ = ~\new_Multi8|ADD16(52)|00_  & ~new_n1718_;
  assign \new_Multi8|x4_01_  = ~new_n1720_ & ~new_n1722_;
  assign \new_Multi8|ADD16(52)|01_  = new_n1714_ | new_n1720_;
  assign new_n1726_ = \new_Multi8|x3_02_  & \new_Multi8|y3_02_ ;
  assign new_n1728_ = ~\new_Multi8|x3_02_  & ~\new_Multi8|y3_02_ ;
  assign new_n1730_ = ~new_n1726_ & ~new_n1728_;
  assign new_n1732_ = \new_Multi8|ADD16(52)|01_  & new_n1730_;
  assign new_n1734_ = ~\new_Multi8|ADD16(52)|01_  & ~new_n1730_;
  assign \new_Multi8|x4_02_  = ~new_n1732_ & ~new_n1734_;
  assign \new_Multi8|ADD16(52)|02_  = new_n1726_ | new_n1732_;
  assign new_n1738_ = \new_Multi8|x3_03_  & \new_Multi8|y3_03_ ;
  assign new_n1740_ = ~\new_Multi8|x3_03_  & ~\new_Multi8|y3_03_ ;
  assign new_n1742_ = ~new_n1738_ & ~new_n1740_;
  assign new_n1744_ = \new_Multi8|ADD16(52)|02_  & new_n1742_;
  assign new_n1746_ = ~\new_Multi8|ADD16(52)|02_  & ~new_n1742_;
  assign \new_Multi8|x4_03_  = ~new_n1744_ & ~new_n1746_;
  assign \new_Multi8|ADD16(52)|03_  = new_n1738_ | new_n1744_;
  assign new_n1750_ = \new_Multi8|x3_04_  & \new_Multi8|y3_04_ ;
  assign new_n1752_ = ~\new_Multi8|x3_04_  & ~\new_Multi8|y3_04_ ;
  assign new_n1754_ = ~new_n1750_ & ~new_n1752_;
  assign new_n1756_ = \new_Multi8|ADD16(52)|03_  & new_n1754_;
  assign new_n1758_ = ~\new_Multi8|ADD16(52)|03_  & ~new_n1754_;
  assign \new_Multi8|x4_04_  = ~new_n1756_ & ~new_n1758_;
  assign \new_Multi8|ADD16(52)|04_  = new_n1750_ | new_n1756_;
  assign new_n1762_ = \new_Multi8|x3_05_  & \new_Multi8|y3_05_ ;
  assign new_n1764_ = ~\new_Multi8|x3_05_  & ~\new_Multi8|y3_05_ ;
  assign new_n1766_ = ~new_n1762_ & ~new_n1764_;
  assign new_n1768_ = \new_Multi8|ADD16(52)|04_  & new_n1766_;
  assign new_n1770_ = ~\new_Multi8|ADD16(52)|04_  & ~new_n1766_;
  assign \new_Multi8|x4_05_  = ~new_n1768_ & ~new_n1770_;
  assign \new_Multi8|ADD16(52)|05_  = new_n1762_ | new_n1768_;
  assign new_n1774_ = \new_Multi8|x3_06_  & \new_Multi8|y3_06_ ;
  assign new_n1776_ = ~\new_Multi8|x3_06_  & ~\new_Multi8|y3_06_ ;
  assign new_n1778_ = ~new_n1774_ & ~new_n1776_;
  assign new_n1780_ = \new_Multi8|ADD16(52)|05_  & new_n1778_;
  assign new_n1782_ = ~\new_Multi8|ADD16(52)|05_  & ~new_n1778_;
  assign \new_Multi8|x4_06_  = ~new_n1780_ & ~new_n1782_;
  assign \new_Multi8|ADD16(52)|06_  = new_n1774_ | new_n1780_;
  assign new_n1786_ = \new_Multi8|x3_07_  & \new_Multi8|y3_07_ ;
  assign new_n1788_ = ~\new_Multi8|x3_07_  & ~\new_Multi8|y3_07_ ;
  assign new_n1790_ = ~new_n1786_ & ~new_n1788_;
  assign new_n1792_ = \new_Multi8|ADD16(52)|06_  & new_n1790_;
  assign new_n1794_ = ~\new_Multi8|ADD16(52)|06_  & ~new_n1790_;
  assign \new_Multi8|x4_07_  = ~new_n1792_ & ~new_n1794_;
  assign \new_Multi8|ADD16(52)|07_  = new_n1786_ | new_n1792_;
  assign new_n1798_ = \new_Multi8|x3_08_  & \new_Multi8|y3_08_ ;
  assign new_n1800_ = ~\new_Multi8|x3_08_  & ~\new_Multi8|y3_08_ ;
  assign new_n1802_ = ~new_n1798_ & ~new_n1800_;
  assign new_n1804_ = \new_Multi8|ADD16(52)|07_  & new_n1802_;
  assign new_n1806_ = ~\new_Multi8|ADD16(52)|07_  & ~new_n1802_;
  assign \new_Multi8|x4_08_  = ~new_n1804_ & ~new_n1806_;
  assign \new_Multi8|ADD16(52)|08_  = new_n1798_ | new_n1804_;
  assign new_n1810_ = \new_Multi8|x3_09_  & \new_Multi8|y3_09_ ;
  assign new_n1812_ = ~\new_Multi8|x3_09_  & ~\new_Multi8|y3_09_ ;
  assign new_n1814_ = ~new_n1810_ & ~new_n1812_;
  assign new_n1816_ = \new_Multi8|ADD16(52)|08_  & new_n1814_;
  assign new_n1818_ = ~\new_Multi8|ADD16(52)|08_  & ~new_n1814_;
  assign \new_Multi8|x4_09_  = ~new_n1816_ & ~new_n1818_;
  assign \new_Multi8|ADD16(52)|09_  = new_n1810_ | new_n1816_;
  assign new_n1822_ = \new_Multi8|x3_10_  & \new_Multi8|y3_10_ ;
  assign new_n1824_ = ~\new_Multi8|x3_10_  & ~\new_Multi8|y3_10_ ;
  assign new_n1826_ = ~new_n1822_ & ~new_n1824_;
  assign new_n1828_ = \new_Multi8|ADD16(52)|09_  & new_n1826_;
  assign new_n1830_ = ~\new_Multi8|ADD16(52)|09_  & ~new_n1826_;
  assign \new_Multi8|x4_10_  = ~new_n1828_ & ~new_n1830_;
  assign \new_Multi8|ADD16(52)|10_  = new_n1822_ | new_n1828_;
  assign new_n1834_ = \new_Multi8|x3_11_  & \new_Multi8|y3_11_ ;
  assign new_n1836_ = ~\new_Multi8|x3_11_  & ~\new_Multi8|y3_11_ ;
  assign new_n1838_ = ~new_n1834_ & ~new_n1836_;
  assign new_n1840_ = \new_Multi8|ADD16(52)|10_  & new_n1838_;
  assign new_n1842_ = ~\new_Multi8|ADD16(52)|10_  & ~new_n1838_;
  assign \new_Multi8|x4_11_  = ~new_n1840_ & ~new_n1842_;
  assign \new_Multi8|ADD16(52)|11_  = new_n1834_ | new_n1840_;
  assign new_n1846_ = \new_Multi8|x3_12_  & \new_Multi8|y3_12_ ;
  assign new_n1848_ = ~\new_Multi8|x3_12_  & ~\new_Multi8|y3_12_ ;
  assign new_n1850_ = ~new_n1846_ & ~new_n1848_;
  assign new_n1852_ = \new_Multi8|ADD16(52)|11_  & new_n1850_;
  assign new_n1854_ = ~\new_Multi8|ADD16(52)|11_  & ~new_n1850_;
  assign \new_Multi8|x4_12_  = ~new_n1852_ & ~new_n1854_;
  assign \new_Multi8|ADD16(52)|12_  = new_n1846_ | new_n1852_;
  assign new_n1858_ = \new_Multi8|x3_13_  & \new_Multi8|y3_13_ ;
  assign new_n1860_ = ~\new_Multi8|x3_13_  & ~\new_Multi8|y3_13_ ;
  assign new_n1862_ = ~new_n1858_ & ~new_n1860_;
  assign new_n1864_ = \new_Multi8|ADD16(52)|12_  & new_n1862_;
  assign new_n1866_ = ~\new_Multi8|ADD16(52)|12_  & ~new_n1862_;
  assign \new_Multi8|x4_13_  = ~new_n1864_ & ~new_n1866_;
  assign \new_Multi8|ADD16(52)|13_  = new_n1858_ | new_n1864_;
  assign new_n1870_ = \new_Multi8|x3_14_  & \new_Multi8|y3_14_ ;
  assign new_n1872_ = ~\new_Multi8|x3_14_  & ~\new_Multi8|y3_14_ ;
  assign new_n1874_ = ~new_n1870_ & ~new_n1872_;
  assign new_n1876_ = \new_Multi8|ADD16(52)|13_  & new_n1874_;
  assign new_n1878_ = ~\new_Multi8|ADD16(52)|13_  & ~new_n1874_;
  assign \new_Multi8|x4_14_  = ~new_n1876_ & ~new_n1878_;
  assign \new_Multi8|ADD16(52)|14_  = new_n1870_ | new_n1876_;
  assign new_n1882_ = \new_Multi8|x3_15_  & \new_Multi8|y3_15_ ;
  assign new_n1884_ = ~\new_Multi8|x3_15_  & ~\new_Multi8|y3_15_ ;
  assign new_n1886_ = ~new_n1882_ & ~new_n1884_;
  assign new_n1888_ = \new_Multi8|ADD16(52)|14_  & new_n1886_;
  assign new_n1890_ = ~\new_Multi8|ADD16(52)|14_  & ~new_n1886_;
  assign \new_Multi8|x4_15_  = ~new_n1888_ & ~new_n1890_;
  assign \new_Multi8|ADD16(69)|c_  = 1'b0;
  assign new_n1911_ = \new_Multi8|x4_00_  & \new_Multi8|y4_00_ ;
  assign new_n1913_ = ~\new_Multi8|x4_00_  & ~\new_Multi8|y4_00_ ;
  assign new_n1915_ = ~new_n1911_ & ~new_n1913_;
  assign new_n1917_ = \new_Multi8|ADD16(69)|c_  & new_n1915_;
  assign new_n1919_ = ~\new_Multi8|ADD16(69)|c_  & ~new_n1915_;
  assign \new_Multi8|x5_00_  = ~new_n1917_ & ~new_n1919_;
  assign \new_Multi8|ADD16(69)|00_  = new_n1911_ | new_n1917_;
  assign new_n1923_ = \new_Multi8|x4_01_  & \new_Multi8|y4_01_ ;
  assign new_n1925_ = ~\new_Multi8|x4_01_  & ~\new_Multi8|y4_01_ ;
  assign new_n1927_ = ~new_n1923_ & ~new_n1925_;
  assign new_n1929_ = \new_Multi8|ADD16(69)|00_  & new_n1927_;
  assign new_n1931_ = ~\new_Multi8|ADD16(69)|00_  & ~new_n1927_;
  assign \new_Multi8|x5_01_  = ~new_n1929_ & ~new_n1931_;
  assign \new_Multi8|ADD16(69)|01_  = new_n1923_ | new_n1929_;
  assign new_n1935_ = \new_Multi8|x4_02_  & \new_Multi8|y4_02_ ;
  assign new_n1937_ = ~\new_Multi8|x4_02_  & ~\new_Multi8|y4_02_ ;
  assign new_n1939_ = ~new_n1935_ & ~new_n1937_;
  assign new_n1941_ = \new_Multi8|ADD16(69)|01_  & new_n1939_;
  assign new_n1943_ = ~\new_Multi8|ADD16(69)|01_  & ~new_n1939_;
  assign \new_Multi8|x5_02_  = ~new_n1941_ & ~new_n1943_;
  assign \new_Multi8|ADD16(69)|02_  = new_n1935_ | new_n1941_;
  assign new_n1947_ = \new_Multi8|x4_03_  & \new_Multi8|y4_03_ ;
  assign new_n1949_ = ~\new_Multi8|x4_03_  & ~\new_Multi8|y4_03_ ;
  assign new_n1951_ = ~new_n1947_ & ~new_n1949_;
  assign new_n1953_ = \new_Multi8|ADD16(69)|02_  & new_n1951_;
  assign new_n1955_ = ~\new_Multi8|ADD16(69)|02_  & ~new_n1951_;
  assign \new_Multi8|x5_03_  = ~new_n1953_ & ~new_n1955_;
  assign \new_Multi8|ADD16(69)|03_  = new_n1947_ | new_n1953_;
  assign new_n1959_ = \new_Multi8|x4_04_  & \new_Multi8|y4_04_ ;
  assign new_n1961_ = ~\new_Multi8|x4_04_  & ~\new_Multi8|y4_04_ ;
  assign new_n1963_ = ~new_n1959_ & ~new_n1961_;
  assign new_n1965_ = \new_Multi8|ADD16(69)|03_  & new_n1963_;
  assign new_n1967_ = ~\new_Multi8|ADD16(69)|03_  & ~new_n1963_;
  assign \new_Multi8|x5_04_  = ~new_n1965_ & ~new_n1967_;
  assign \new_Multi8|ADD16(69)|04_  = new_n1959_ | new_n1965_;
  assign new_n1971_ = \new_Multi8|x4_05_  & \new_Multi8|y4_05_ ;
  assign new_n1973_ = ~\new_Multi8|x4_05_  & ~\new_Multi8|y4_05_ ;
  assign new_n1975_ = ~new_n1971_ & ~new_n1973_;
  assign new_n1977_ = \new_Multi8|ADD16(69)|04_  & new_n1975_;
  assign new_n1979_ = ~\new_Multi8|ADD16(69)|04_  & ~new_n1975_;
  assign \new_Multi8|x5_05_  = ~new_n1977_ & ~new_n1979_;
  assign \new_Multi8|ADD16(69)|05_  = new_n1971_ | new_n1977_;
  assign new_n1983_ = \new_Multi8|x4_06_  & \new_Multi8|y4_06_ ;
  assign new_n1985_ = ~\new_Multi8|x4_06_  & ~\new_Multi8|y4_06_ ;
  assign new_n1987_ = ~new_n1983_ & ~new_n1985_;
  assign new_n1989_ = \new_Multi8|ADD16(69)|05_  & new_n1987_;
  assign new_n1991_ = ~\new_Multi8|ADD16(69)|05_  & ~new_n1987_;
  assign \new_Multi8|x5_06_  = ~new_n1989_ & ~new_n1991_;
  assign \new_Multi8|ADD16(69)|06_  = new_n1983_ | new_n1989_;
  assign new_n1995_ = \new_Multi8|x4_07_  & \new_Multi8|y4_07_ ;
  assign new_n1997_ = ~\new_Multi8|x4_07_  & ~\new_Multi8|y4_07_ ;
  assign new_n1999_ = ~new_n1995_ & ~new_n1997_;
  assign new_n2001_ = \new_Multi8|ADD16(69)|06_  & new_n1999_;
  assign new_n2003_ = ~\new_Multi8|ADD16(69)|06_  & ~new_n1999_;
  assign \new_Multi8|x5_07_  = ~new_n2001_ & ~new_n2003_;
  assign \new_Multi8|ADD16(69)|07_  = new_n1995_ | new_n2001_;
  assign new_n2007_ = \new_Multi8|x4_08_  & \new_Multi8|y4_08_ ;
  assign new_n2009_ = ~\new_Multi8|x4_08_  & ~\new_Multi8|y4_08_ ;
  assign new_n2011_ = ~new_n2007_ & ~new_n2009_;
  assign new_n2013_ = \new_Multi8|ADD16(69)|07_  & new_n2011_;
  assign new_n2015_ = ~\new_Multi8|ADD16(69)|07_  & ~new_n2011_;
  assign \new_Multi8|x5_08_  = ~new_n2013_ & ~new_n2015_;
  assign \new_Multi8|ADD16(69)|08_  = new_n2007_ | new_n2013_;
  assign new_n2019_ = \new_Multi8|x4_09_  & \new_Multi8|y4_09_ ;
  assign new_n2021_ = ~\new_Multi8|x4_09_  & ~\new_Multi8|y4_09_ ;
  assign new_n2023_ = ~new_n2019_ & ~new_n2021_;
  assign new_n2025_ = \new_Multi8|ADD16(69)|08_  & new_n2023_;
  assign new_n2027_ = ~\new_Multi8|ADD16(69)|08_  & ~new_n2023_;
  assign \new_Multi8|x5_09_  = ~new_n2025_ & ~new_n2027_;
  assign \new_Multi8|ADD16(69)|09_  = new_n2019_ | new_n2025_;
  assign new_n2031_ = \new_Multi8|x4_10_  & \new_Multi8|y4_10_ ;
  assign new_n2033_ = ~\new_Multi8|x4_10_  & ~\new_Multi8|y4_10_ ;
  assign new_n2035_ = ~new_n2031_ & ~new_n2033_;
  assign new_n2037_ = \new_Multi8|ADD16(69)|09_  & new_n2035_;
  assign new_n2039_ = ~\new_Multi8|ADD16(69)|09_  & ~new_n2035_;
  assign \new_Multi8|x5_10_  = ~new_n2037_ & ~new_n2039_;
  assign \new_Multi8|ADD16(69)|10_  = new_n2031_ | new_n2037_;
  assign new_n2043_ = \new_Multi8|x4_11_  & \new_Multi8|y4_11_ ;
  assign new_n2045_ = ~\new_Multi8|x4_11_  & ~\new_Multi8|y4_11_ ;
  assign new_n2047_ = ~new_n2043_ & ~new_n2045_;
  assign new_n2049_ = \new_Multi8|ADD16(69)|10_  & new_n2047_;
  assign new_n2051_ = ~\new_Multi8|ADD16(69)|10_  & ~new_n2047_;
  assign \new_Multi8|x5_11_  = ~new_n2049_ & ~new_n2051_;
  assign \new_Multi8|ADD16(69)|11_  = new_n2043_ | new_n2049_;
  assign new_n2055_ = \new_Multi8|x4_12_  & \new_Multi8|y4_12_ ;
  assign new_n2057_ = ~\new_Multi8|x4_12_  & ~\new_Multi8|y4_12_ ;
  assign new_n2059_ = ~new_n2055_ & ~new_n2057_;
  assign new_n2061_ = \new_Multi8|ADD16(69)|11_  & new_n2059_;
  assign new_n2063_ = ~\new_Multi8|ADD16(69)|11_  & ~new_n2059_;
  assign \new_Multi8|x5_12_  = ~new_n2061_ & ~new_n2063_;
  assign \new_Multi8|ADD16(69)|12_  = new_n2055_ | new_n2061_;
  assign new_n2067_ = \new_Multi8|x4_13_  & \new_Multi8|y4_13_ ;
  assign new_n2069_ = ~\new_Multi8|x4_13_  & ~\new_Multi8|y4_13_ ;
  assign new_n2071_ = ~new_n2067_ & ~new_n2069_;
  assign new_n2073_ = \new_Multi8|ADD16(69)|12_  & new_n2071_;
  assign new_n2075_ = ~\new_Multi8|ADD16(69)|12_  & ~new_n2071_;
  assign \new_Multi8|x5_13_  = ~new_n2073_ & ~new_n2075_;
  assign \new_Multi8|ADD16(69)|13_  = new_n2067_ | new_n2073_;
  assign new_n2079_ = \new_Multi8|x4_14_  & \new_Multi8|y4_14_ ;
  assign new_n2081_ = ~\new_Multi8|x4_14_  & ~\new_Multi8|y4_14_ ;
  assign new_n2083_ = ~new_n2079_ & ~new_n2081_;
  assign new_n2085_ = \new_Multi8|ADD16(69)|13_  & new_n2083_;
  assign new_n2087_ = ~\new_Multi8|ADD16(69)|13_  & ~new_n2083_;
  assign \new_Multi8|x5_14_  = ~new_n2085_ & ~new_n2087_;
  assign \new_Multi8|ADD16(69)|14_  = new_n2079_ | new_n2085_;
  assign new_n2091_ = \new_Multi8|x4_15_  & \new_Multi8|y4_15_ ;
  assign new_n2093_ = ~\new_Multi8|x4_15_  & ~\new_Multi8|y4_15_ ;
  assign new_n2095_ = ~new_n2091_ & ~new_n2093_;
  assign new_n2097_ = \new_Multi8|ADD16(69)|14_  & new_n2095_;
  assign new_n2099_ = ~\new_Multi8|ADD16(69)|14_  & ~new_n2095_;
  assign \new_Multi8|x5_15_  = ~new_n2097_ & ~new_n2099_;
endmodule


