// Benchmark "ADD100" written by ABC on Tue Apr  9 09:11:33 2024

module ADD100 ( 
    a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a10, a11, a12, a13,
    a14, a15, a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27,
    a28, a29, a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40, a41,
    a42, a43, a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54, a55,
    a56, a57, a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68, a69,
    a70, a71, a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82, a83,
    a84, a85, a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96, a97,
    a98, a99, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b10, b11,
    b12, b13, b14, b15, b16, b17, b18, b19, b20, b21, b22, b23, b24, b25,
    b26, b27, b28, b29, b30, b31, b32, b33, b34, b35, b36, b37, b38, b39,
    b40, b41, b42, b43, b44, b45, b46, b47, b48, b49, b50, b51, b52, b53,
    b54, b55, b56, b57, b58, b59, b60, b61, b62, b63, b64, b65, b66, b67,
    b68, b69, b70, b71, b72, b73, b74, b75, b76, b77, b78, b79, b80, b81,
    b82, b83, b84, b85, b86, b87, b88, b89, b90, b91, b92, b93, b94, b95,
    b96, b97, b98, b99,
    s00, s01, s02, s03, s04, s05, s06, s07, s08, s09, s10, s11, s12, s13,
    s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27,
    s28, s29, s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41,
    s42, s43, s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55,
    s56, s57, s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69,
    s70, s71, s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83,
    s84, s85, s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97,
    s98, s99, s100  );
  input  a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a10, a11, a12,
    a13, a14, a15, a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26,
    a27, a28, a29, a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40,
    a41, a42, a43, a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54,
    a55, a56, a57, a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68,
    a69, a70, a71, a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82,
    a83, a84, a85, a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96,
    a97, a98, a99, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b10,
    b11, b12, b13, b14, b15, b16, b17, b18, b19, b20, b21, b22, b23, b24,
    b25, b26, b27, b28, b29, b30, b31, b32, b33, b34, b35, b36, b37, b38,
    b39, b40, b41, b42, b43, b44, b45, b46, b47, b48, b49, b50, b51, b52,
    b53, b54, b55, b56, b57, b58, b59, b60, b61, b62, b63, b64, b65, b66,
    b67, b68, b69, b70, b71, b72, b73, b74, b75, b76, b77, b78, b79, b80,
    b81, b82, b83, b84, b85, b86, b87, b88, b89, b90, b91, b92, b93, b94,
    b95, b96, b97, b98, b99;
  output s00, s01, s02, s03, s04, s05, s06, s07, s08, s09, s10, s11, s12, s13,
    s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27,
    s28, s29, s30, s31, s32, s33, s34, s35, s36, s37, s38, s39, s40, s41,
    s42, s43, s44, s45, s46, s47, s48, s49, s50, s51, s52, s53, s54, s55,
    s56, s57, s58, s59, s60, s61, s62, s63, s64, s65, s66, s67, s68, s69,
    s70, s71, s72, s73, s74, s75, s76, s77, s78, s79, s80, s81, s82, s83,
    s84, s85, s86, s87, s88, s89, s90, s91, s92, s93, s94, s95, s96, s97,
    s98, s99, s100;
  wire \new_ADD100|c_ , new_n704_, new_n706_, new_n708_, new_n710_,
    new_n712_, \new_ADD100|00_ , new_n716_, new_n718_, new_n720_,
    new_n722_, new_n724_, \new_ADD100|01_ , new_n728_, new_n730_,
    new_n732_, new_n734_, new_n736_, \new_ADD100|02_ , new_n740_,
    new_n742_, new_n744_, new_n746_, new_n748_, \new_ADD100|03_ ,
    new_n752_, new_n754_, new_n756_, new_n758_, new_n760_,
    \new_ADD100|04_ , new_n764_, new_n766_, new_n768_, new_n770_,
    new_n772_, \new_ADD100|05_ , new_n776_, new_n778_, new_n780_,
    new_n782_, new_n784_, \new_ADD100|06_ , new_n788_, new_n790_,
    new_n792_, new_n794_, new_n796_, \new_ADD100|07_ , new_n800_,
    new_n802_, new_n804_, new_n806_, new_n808_, \new_ADD100|08_ ,
    new_n812_, new_n814_, new_n816_, new_n818_, new_n820_,
    \new_ADD100|09_ , new_n824_, new_n826_, new_n828_, new_n830_,
    new_n832_, \new_ADD100|10_ , new_n836_, new_n838_, new_n840_,
    new_n842_, new_n844_, \new_ADD100|11_ , new_n848_, new_n850_,
    new_n852_, new_n854_, new_n856_, \new_ADD100|12_ , new_n860_,
    new_n862_, new_n864_, new_n866_, new_n868_, \new_ADD100|13_ ,
    new_n872_, new_n874_, new_n876_, new_n878_, new_n880_,
    \new_ADD100|14_ , new_n884_, new_n886_, new_n888_, new_n890_,
    new_n892_, \new_ADD100|15_ , new_n896_, new_n898_, new_n900_,
    new_n902_, new_n904_, \new_ADD100|16_ , new_n908_, new_n910_,
    new_n912_, new_n914_, new_n916_, \new_ADD100|17_ , new_n920_,
    new_n922_, new_n924_, new_n926_, new_n928_, \new_ADD100|18_ ,
    new_n932_, new_n934_, new_n936_, new_n938_, new_n940_,
    \new_ADD100|19_ , new_n944_, new_n946_, new_n948_, new_n950_,
    new_n952_, \new_ADD100|20_ , new_n956_, new_n958_, new_n960_,
    new_n962_, new_n964_, \new_ADD100|21_ , new_n968_, new_n970_,
    new_n972_, new_n974_, new_n976_, \new_ADD100|22_ , new_n980_,
    new_n982_, new_n984_, new_n986_, new_n988_, \new_ADD100|23_ ,
    new_n992_, new_n994_, new_n996_, new_n998_, new_n1000_,
    \new_ADD100|24_ , new_n1004_, new_n1006_, new_n1008_, new_n1010_,
    new_n1012_, \new_ADD100|25_ , new_n1016_, new_n1018_, new_n1020_,
    new_n1022_, new_n1024_, \new_ADD100|26_ , new_n1028_, new_n1030_,
    new_n1032_, new_n1034_, new_n1036_, \new_ADD100|27_ , new_n1040_,
    new_n1042_, new_n1044_, new_n1046_, new_n1048_, \new_ADD100|28_ ,
    new_n1052_, new_n1054_, new_n1056_, new_n1058_, new_n1060_,
    \new_ADD100|29_ , new_n1064_, new_n1066_, new_n1068_, new_n1070_,
    new_n1072_, \new_ADD100|30_ , new_n1076_, new_n1078_, new_n1080_,
    new_n1082_, new_n1084_, \new_ADD100|31_ , new_n1088_, new_n1090_,
    new_n1092_, new_n1094_, new_n1096_, \new_ADD100|32_ , new_n1100_,
    new_n1102_, new_n1104_, new_n1106_, new_n1108_, \new_ADD100|33_ ,
    new_n1112_, new_n1114_, new_n1116_, new_n1118_, new_n1120_,
    \new_ADD100|34_ , new_n1124_, new_n1126_, new_n1128_, new_n1130_,
    new_n1132_, \new_ADD100|35_ , new_n1136_, new_n1138_, new_n1140_,
    new_n1142_, new_n1144_, \new_ADD100|36_ , new_n1148_, new_n1150_,
    new_n1152_, new_n1154_, new_n1156_, \new_ADD100|37_ , new_n1160_,
    new_n1162_, new_n1164_, new_n1166_, new_n1168_, \new_ADD100|38_ ,
    new_n1172_, new_n1174_, new_n1176_, new_n1178_, new_n1180_,
    \new_ADD100|39_ , new_n1184_, new_n1186_, new_n1188_, new_n1190_,
    new_n1192_, \new_ADD100|40_ , new_n1196_, new_n1198_, new_n1200_,
    new_n1202_, new_n1204_, \new_ADD100|41_ , new_n1208_, new_n1210_,
    new_n1212_, new_n1214_, new_n1216_, \new_ADD100|42_ , new_n1220_,
    new_n1222_, new_n1224_, new_n1226_, new_n1228_, \new_ADD100|43_ ,
    new_n1232_, new_n1234_, new_n1236_, new_n1238_, new_n1240_,
    \new_ADD100|44_ , new_n1244_, new_n1246_, new_n1248_, new_n1250_,
    new_n1252_, \new_ADD100|45_ , new_n1256_, new_n1258_, new_n1260_,
    new_n1262_, new_n1264_, \new_ADD100|46_ , new_n1268_, new_n1270_,
    new_n1272_, new_n1274_, new_n1276_, \new_ADD100|47_ , new_n1280_,
    new_n1282_, new_n1284_, new_n1286_, new_n1288_, \new_ADD100|48_ ,
    new_n1292_, new_n1294_, new_n1296_, new_n1298_, new_n1300_,
    \new_ADD100|49_ , new_n1304_, new_n1306_, new_n1308_, new_n1310_,
    new_n1312_, \new_ADD100|50_ , new_n1316_, new_n1318_, new_n1320_,
    new_n1322_, new_n1324_, \new_ADD100|51_ , new_n1328_, new_n1330_,
    new_n1332_, new_n1334_, new_n1336_, \new_ADD100|52_ , new_n1340_,
    new_n1342_, new_n1344_, new_n1346_, new_n1348_, \new_ADD100|53_ ,
    new_n1352_, new_n1354_, new_n1356_, new_n1358_, new_n1360_,
    \new_ADD100|54_ , new_n1364_, new_n1366_, new_n1368_, new_n1370_,
    new_n1372_, \new_ADD100|55_ , new_n1376_, new_n1378_, new_n1380_,
    new_n1382_, new_n1384_, \new_ADD100|56_ , new_n1388_, new_n1390_,
    new_n1392_, new_n1394_, new_n1396_, \new_ADD100|57_ , new_n1400_,
    new_n1402_, new_n1404_, new_n1406_, new_n1408_, \new_ADD100|58_ ,
    new_n1412_, new_n1414_, new_n1416_, new_n1418_, new_n1420_,
    \new_ADD100|59_ , new_n1424_, new_n1426_, new_n1428_, new_n1430_,
    new_n1432_, \new_ADD100|60_ , new_n1436_, new_n1438_, new_n1440_,
    new_n1442_, new_n1444_, \new_ADD100|61_ , new_n1448_, new_n1450_,
    new_n1452_, new_n1454_, new_n1456_, \new_ADD100|62_ , new_n1460_,
    new_n1462_, new_n1464_, new_n1466_, new_n1468_, \new_ADD100|63_ ,
    new_n1472_, new_n1474_, new_n1476_, new_n1478_, new_n1480_,
    \new_ADD100|64_ , new_n1484_, new_n1486_, new_n1488_, new_n1490_,
    new_n1492_, \new_ADD100|65_ , new_n1496_, new_n1498_, new_n1500_,
    new_n1502_, new_n1504_, \new_ADD100|66_ , new_n1508_, new_n1510_,
    new_n1512_, new_n1514_, new_n1516_, \new_ADD100|67_ , new_n1520_,
    new_n1522_, new_n1524_, new_n1526_, new_n1528_, \new_ADD100|68_ ,
    new_n1532_, new_n1534_, new_n1536_, new_n1538_, new_n1540_,
    \new_ADD100|69_ , new_n1544_, new_n1546_, new_n1548_, new_n1550_,
    new_n1552_, \new_ADD100|70_ , new_n1556_, new_n1558_, new_n1560_,
    new_n1562_, new_n1564_, \new_ADD100|71_ , new_n1568_, new_n1570_,
    new_n1572_, new_n1574_, new_n1576_, \new_ADD100|72_ , new_n1580_,
    new_n1582_, new_n1584_, new_n1586_, new_n1588_, \new_ADD100|73_ ,
    new_n1592_, new_n1594_, new_n1596_, new_n1598_, new_n1600_,
    \new_ADD100|74_ , new_n1604_, new_n1606_, new_n1608_, new_n1610_,
    new_n1612_, \new_ADD100|75_ , new_n1616_, new_n1618_, new_n1620_,
    new_n1622_, new_n1624_, \new_ADD100|76_ , new_n1628_, new_n1630_,
    new_n1632_, new_n1634_, new_n1636_, \new_ADD100|77_ , new_n1640_,
    new_n1642_, new_n1644_, new_n1646_, new_n1648_, \new_ADD100|78_ ,
    new_n1652_, new_n1654_, new_n1656_, new_n1658_, new_n1660_,
    \new_ADD100|79_ , new_n1664_, new_n1666_, new_n1668_, new_n1670_,
    new_n1672_, \new_ADD100|80_ , new_n1676_, new_n1678_, new_n1680_,
    new_n1682_, new_n1684_, \new_ADD100|81_ , new_n1688_, new_n1690_,
    new_n1692_, new_n1694_, new_n1696_, \new_ADD100|82_ , new_n1700_,
    new_n1702_, new_n1704_, new_n1706_, new_n1708_, \new_ADD100|83_ ,
    new_n1712_, new_n1714_, new_n1716_, new_n1718_, new_n1720_,
    \new_ADD100|84_ , new_n1724_, new_n1726_, new_n1728_, new_n1730_,
    new_n1732_, \new_ADD100|85_ , new_n1736_, new_n1738_, new_n1740_,
    new_n1742_, new_n1744_, \new_ADD100|86_ , new_n1748_, new_n1750_,
    new_n1752_, new_n1754_, new_n1756_, \new_ADD100|87_ , new_n1760_,
    new_n1762_, new_n1764_, new_n1766_, new_n1768_, \new_ADD100|88_ ,
    new_n1772_, new_n1774_, new_n1776_, new_n1778_, new_n1780_,
    \new_ADD100|89_ , new_n1784_, new_n1786_, new_n1788_, new_n1790_,
    new_n1792_, \new_ADD100|90_ , new_n1796_, new_n1798_, new_n1800_,
    new_n1802_, new_n1804_, \new_ADD100|91_ , new_n1808_, new_n1810_,
    new_n1812_, new_n1814_, new_n1816_, \new_ADD100|92_ , new_n1820_,
    new_n1822_, new_n1824_, new_n1826_, new_n1828_, \new_ADD100|93_ ,
    new_n1832_, new_n1834_, new_n1836_, new_n1838_, new_n1840_,
    \new_ADD100|94_ , new_n1844_, new_n1846_, new_n1848_, new_n1850_,
    new_n1852_, \new_ADD100|95_ , new_n1856_, new_n1858_, new_n1860_,
    new_n1862_, new_n1864_, \new_ADD100|96_ , new_n1868_, new_n1870_,
    new_n1872_, new_n1874_, new_n1876_, \new_ADD100|97_ , new_n1880_,
    new_n1882_, new_n1884_, new_n1886_, new_n1888_, \new_ADD100|98_ ,
    new_n1892_, new_n1894_, new_n1896_, new_n1898_, new_n1900_;
  assign \new_ADD100|c_  = 1'b0;
  assign new_n704_ = a00 & b00;
  assign new_n706_ = ~a00 & ~b00;
  assign new_n708_ = ~new_n704_ & ~new_n706_;
  assign new_n710_ = \new_ADD100|c_  & new_n708_;
  assign new_n712_ = ~\new_ADD100|c_  & ~new_n708_;
  assign s00 = ~new_n710_ & ~new_n712_;
  assign \new_ADD100|00_  = new_n704_ | new_n710_;
  assign new_n716_ = a01 & b01;
  assign new_n718_ = ~a01 & ~b01;
  assign new_n720_ = ~new_n716_ & ~new_n718_;
  assign new_n722_ = \new_ADD100|00_  & new_n720_;
  assign new_n724_ = ~\new_ADD100|00_  & ~new_n720_;
  assign s01 = ~new_n722_ & ~new_n724_;
  assign \new_ADD100|01_  = new_n716_ | new_n722_;
  assign new_n728_ = a02 & b02;
  assign new_n730_ = ~a02 & ~b02;
  assign new_n732_ = ~new_n728_ & ~new_n730_;
  assign new_n734_ = \new_ADD100|01_  & new_n732_;
  assign new_n736_ = ~\new_ADD100|01_  & ~new_n732_;
  assign s02 = ~new_n734_ & ~new_n736_;
  assign \new_ADD100|02_  = new_n728_ | new_n734_;
  assign new_n740_ = a03 & b03;
  assign new_n742_ = ~a03 & ~b03;
  assign new_n744_ = ~new_n740_ & ~new_n742_;
  assign new_n746_ = \new_ADD100|02_  & new_n744_;
  assign new_n748_ = ~\new_ADD100|02_  & ~new_n744_;
  assign s03 = ~new_n746_ & ~new_n748_;
  assign \new_ADD100|03_  = new_n740_ | new_n746_;
  assign new_n752_ = a04 & b04;
  assign new_n754_ = ~a04 & ~b04;
  assign new_n756_ = ~new_n752_ & ~new_n754_;
  assign new_n758_ = \new_ADD100|03_  & new_n756_;
  assign new_n760_ = ~\new_ADD100|03_  & ~new_n756_;
  assign s04 = ~new_n758_ & ~new_n760_;
  assign \new_ADD100|04_  = new_n752_ | new_n758_;
  assign new_n764_ = a05 & b05;
  assign new_n766_ = ~a05 & ~b05;
  assign new_n768_ = ~new_n764_ & ~new_n766_;
  assign new_n770_ = \new_ADD100|04_  & new_n768_;
  assign new_n772_ = ~\new_ADD100|04_  & ~new_n768_;
  assign s05 = ~new_n770_ & ~new_n772_;
  assign \new_ADD100|05_  = new_n764_ | new_n770_;
  assign new_n776_ = a06 & b06;
  assign new_n778_ = ~a06 & ~b06;
  assign new_n780_ = ~new_n776_ & ~new_n778_;
  assign new_n782_ = \new_ADD100|05_  & new_n780_;
  assign new_n784_ = ~\new_ADD100|05_  & ~new_n780_;
  assign s06 = ~new_n782_ & ~new_n784_;
  assign \new_ADD100|06_  = new_n776_ | new_n782_;
  assign new_n788_ = a07 & b07;
  assign new_n790_ = ~a07 & ~b07;
  assign new_n792_ = ~new_n788_ & ~new_n790_;
  assign new_n794_ = \new_ADD100|06_  & new_n792_;
  assign new_n796_ = ~\new_ADD100|06_  & ~new_n792_;
  assign s07 = ~new_n794_ & ~new_n796_;
  assign \new_ADD100|07_  = new_n788_ | new_n794_;
  assign new_n800_ = a08 & b08;
  assign new_n802_ = ~a08 & ~b08;
  assign new_n804_ = ~new_n800_ & ~new_n802_;
  assign new_n806_ = \new_ADD100|07_  & new_n804_;
  assign new_n808_ = ~\new_ADD100|07_  & ~new_n804_;
  assign s08 = ~new_n806_ & ~new_n808_;
  assign \new_ADD100|08_  = new_n800_ | new_n806_;
  assign new_n812_ = a09 & b09;
  assign new_n814_ = ~a09 & ~b09;
  assign new_n816_ = ~new_n812_ & ~new_n814_;
  assign new_n818_ = \new_ADD100|08_  & new_n816_;
  assign new_n820_ = ~\new_ADD100|08_  & ~new_n816_;
  assign s09 = ~new_n818_ & ~new_n820_;
  assign \new_ADD100|09_  = new_n812_ | new_n818_;
  assign new_n824_ = a10 & b10;
  assign new_n826_ = ~a10 & ~b10;
  assign new_n828_ = ~new_n824_ & ~new_n826_;
  assign new_n830_ = \new_ADD100|09_  & new_n828_;
  assign new_n832_ = ~\new_ADD100|09_  & ~new_n828_;
  assign s10 = ~new_n830_ & ~new_n832_;
  assign \new_ADD100|10_  = new_n824_ | new_n830_;
  assign new_n836_ = a11 & b11;
  assign new_n838_ = ~a11 & ~b11;
  assign new_n840_ = ~new_n836_ & ~new_n838_;
  assign new_n842_ = \new_ADD100|10_  & new_n840_;
  assign new_n844_ = ~\new_ADD100|10_  & ~new_n840_;
  assign s11 = ~new_n842_ & ~new_n844_;
  assign \new_ADD100|11_  = new_n836_ | new_n842_;
  assign new_n848_ = a12 & b12;
  assign new_n850_ = ~a12 & ~b12;
  assign new_n852_ = ~new_n848_ & ~new_n850_;
  assign new_n854_ = \new_ADD100|11_  & new_n852_;
  assign new_n856_ = ~\new_ADD100|11_  & ~new_n852_;
  assign s12 = ~new_n854_ & ~new_n856_;
  assign \new_ADD100|12_  = new_n848_ | new_n854_;
  assign new_n860_ = a13 & b13;
  assign new_n862_ = ~a13 & ~b13;
  assign new_n864_ = ~new_n860_ & ~new_n862_;
  assign new_n866_ = \new_ADD100|12_  & new_n864_;
  assign new_n868_ = ~\new_ADD100|12_  & ~new_n864_;
  assign s13 = ~new_n866_ & ~new_n868_;
  assign \new_ADD100|13_  = new_n860_ | new_n866_;
  assign new_n872_ = a14 & b14;
  assign new_n874_ = ~a14 & ~b14;
  assign new_n876_ = ~new_n872_ & ~new_n874_;
  assign new_n878_ = \new_ADD100|13_  & new_n876_;
  assign new_n880_ = ~\new_ADD100|13_  & ~new_n876_;
  assign s14 = ~new_n878_ & ~new_n880_;
  assign \new_ADD100|14_  = new_n872_ | new_n878_;
  assign new_n884_ = a15 & b15;
  assign new_n886_ = ~a15 & ~b15;
  assign new_n888_ = ~new_n884_ & ~new_n886_;
  assign new_n890_ = \new_ADD100|14_  & new_n888_;
  assign new_n892_ = ~\new_ADD100|14_  & ~new_n888_;
  assign s15 = ~new_n890_ & ~new_n892_;
  assign \new_ADD100|15_  = new_n884_ | new_n890_;
  assign new_n896_ = a16 & b16;
  assign new_n898_ = ~a16 & ~b16;
  assign new_n900_ = ~new_n896_ & ~new_n898_;
  assign new_n902_ = \new_ADD100|15_  & new_n900_;
  assign new_n904_ = ~\new_ADD100|15_  & ~new_n900_;
  assign s16 = ~new_n902_ & ~new_n904_;
  assign \new_ADD100|16_  = new_n896_ | new_n902_;
  assign new_n908_ = a17 & b17;
  assign new_n910_ = ~a17 & ~b17;
  assign new_n912_ = ~new_n908_ & ~new_n910_;
  assign new_n914_ = \new_ADD100|16_  & new_n912_;
  assign new_n916_ = ~\new_ADD100|16_  & ~new_n912_;
  assign s17 = ~new_n914_ & ~new_n916_;
  assign \new_ADD100|17_  = new_n908_ | new_n914_;
  assign new_n920_ = a18 & b18;
  assign new_n922_ = ~a18 & ~b18;
  assign new_n924_ = ~new_n920_ & ~new_n922_;
  assign new_n926_ = \new_ADD100|17_  & new_n924_;
  assign new_n928_ = ~\new_ADD100|17_  & ~new_n924_;
  assign s18 = ~new_n926_ & ~new_n928_;
  assign \new_ADD100|18_  = new_n920_ | new_n926_;
  assign new_n932_ = a19 & b19;
  assign new_n934_ = ~a19 & ~b19;
  assign new_n936_ = ~new_n932_ & ~new_n934_;
  assign new_n938_ = \new_ADD100|18_  & new_n936_;
  assign new_n940_ = ~\new_ADD100|18_  & ~new_n936_;
  assign s19 = ~new_n938_ & ~new_n940_;
  assign \new_ADD100|19_  = new_n932_ | new_n938_;
  assign new_n944_ = a20 & b20;
  assign new_n946_ = ~a20 & ~b20;
  assign new_n948_ = ~new_n944_ & ~new_n946_;
  assign new_n950_ = \new_ADD100|19_  & new_n948_;
  assign new_n952_ = ~\new_ADD100|19_  & ~new_n948_;
  assign s20 = ~new_n950_ & ~new_n952_;
  assign \new_ADD100|20_  = new_n944_ | new_n950_;
  assign new_n956_ = a21 & b21;
  assign new_n958_ = ~a21 & ~b21;
  assign new_n960_ = ~new_n956_ & ~new_n958_;
  assign new_n962_ = \new_ADD100|20_  & new_n960_;
  assign new_n964_ = ~\new_ADD100|20_  & ~new_n960_;
  assign s21 = ~new_n962_ & ~new_n964_;
  assign \new_ADD100|21_  = new_n956_ | new_n962_;
  assign new_n968_ = a22 & b22;
  assign new_n970_ = ~a22 & ~b22;
  assign new_n972_ = ~new_n968_ & ~new_n970_;
  assign new_n974_ = \new_ADD100|21_  & new_n972_;
  assign new_n976_ = ~\new_ADD100|21_  & ~new_n972_;
  assign s22 = ~new_n974_ & ~new_n976_;
  assign \new_ADD100|22_  = new_n968_ | new_n974_;
  assign new_n980_ = a23 & b23;
  assign new_n982_ = ~a23 & ~b23;
  assign new_n984_ = ~new_n980_ & ~new_n982_;
  assign new_n986_ = \new_ADD100|22_  & new_n984_;
  assign new_n988_ = ~\new_ADD100|22_  & ~new_n984_;
  assign s23 = ~new_n986_ & ~new_n988_;
  assign \new_ADD100|23_  = new_n980_ | new_n986_;
  assign new_n992_ = a24 & b24;
  assign new_n994_ = ~a24 & ~b24;
  assign new_n996_ = ~new_n992_ & ~new_n994_;
  assign new_n998_ = \new_ADD100|23_  & new_n996_;
  assign new_n1000_ = ~\new_ADD100|23_  & ~new_n996_;
  assign s24 = ~new_n998_ & ~new_n1000_;
  assign \new_ADD100|24_  = new_n992_ | new_n998_;
  assign new_n1004_ = a25 & b25;
  assign new_n1006_ = ~a25 & ~b25;
  assign new_n1008_ = ~new_n1004_ & ~new_n1006_;
  assign new_n1010_ = \new_ADD100|24_  & new_n1008_;
  assign new_n1012_ = ~\new_ADD100|24_  & ~new_n1008_;
  assign s25 = ~new_n1010_ & ~new_n1012_;
  assign \new_ADD100|25_  = new_n1004_ | new_n1010_;
  assign new_n1016_ = a26 & b26;
  assign new_n1018_ = ~a26 & ~b26;
  assign new_n1020_ = ~new_n1016_ & ~new_n1018_;
  assign new_n1022_ = \new_ADD100|25_  & new_n1020_;
  assign new_n1024_ = ~\new_ADD100|25_  & ~new_n1020_;
  assign s26 = ~new_n1022_ & ~new_n1024_;
  assign \new_ADD100|26_  = new_n1016_ | new_n1022_;
  assign new_n1028_ = a27 & b27;
  assign new_n1030_ = ~a27 & ~b27;
  assign new_n1032_ = ~new_n1028_ & ~new_n1030_;
  assign new_n1034_ = \new_ADD100|26_  & new_n1032_;
  assign new_n1036_ = ~\new_ADD100|26_  & ~new_n1032_;
  assign s27 = ~new_n1034_ & ~new_n1036_;
  assign \new_ADD100|27_  = new_n1028_ | new_n1034_;
  assign new_n1040_ = a28 & b28;
  assign new_n1042_ = ~a28 & ~b28;
  assign new_n1044_ = ~new_n1040_ & ~new_n1042_;
  assign new_n1046_ = \new_ADD100|27_  & new_n1044_;
  assign new_n1048_ = ~\new_ADD100|27_  & ~new_n1044_;
  assign s28 = ~new_n1046_ & ~new_n1048_;
  assign \new_ADD100|28_  = new_n1040_ | new_n1046_;
  assign new_n1052_ = a29 & b29;
  assign new_n1054_ = ~a29 & ~b29;
  assign new_n1056_ = ~new_n1052_ & ~new_n1054_;
  assign new_n1058_ = \new_ADD100|28_  & new_n1056_;
  assign new_n1060_ = ~\new_ADD100|28_  & ~new_n1056_;
  assign s29 = ~new_n1058_ & ~new_n1060_;
  assign \new_ADD100|29_  = new_n1052_ | new_n1058_;
  assign new_n1064_ = a30 & b30;
  assign new_n1066_ = ~a30 & ~b30;
  assign new_n1068_ = ~new_n1064_ & ~new_n1066_;
  assign new_n1070_ = \new_ADD100|29_  & new_n1068_;
  assign new_n1072_ = ~\new_ADD100|29_  & ~new_n1068_;
  assign s30 = ~new_n1070_ & ~new_n1072_;
  assign \new_ADD100|30_  = new_n1064_ | new_n1070_;
  assign new_n1076_ = a31 & b31;
  assign new_n1078_ = ~a31 & ~b31;
  assign new_n1080_ = ~new_n1076_ & ~new_n1078_;
  assign new_n1082_ = \new_ADD100|30_  & new_n1080_;
  assign new_n1084_ = ~\new_ADD100|30_  & ~new_n1080_;
  assign s31 = ~new_n1082_ & ~new_n1084_;
  assign \new_ADD100|31_  = new_n1076_ | new_n1082_;
  assign new_n1088_ = a32 & b32;
  assign new_n1090_ = ~a32 & ~b32;
  assign new_n1092_ = ~new_n1088_ & ~new_n1090_;
  assign new_n1094_ = \new_ADD100|31_  & new_n1092_;
  assign new_n1096_ = ~\new_ADD100|31_  & ~new_n1092_;
  assign s32 = ~new_n1094_ & ~new_n1096_;
  assign \new_ADD100|32_  = new_n1088_ | new_n1094_;
  assign new_n1100_ = a33 & b33;
  assign new_n1102_ = ~a33 & ~b33;
  assign new_n1104_ = ~new_n1100_ & ~new_n1102_;
  assign new_n1106_ = \new_ADD100|32_  & new_n1104_;
  assign new_n1108_ = ~\new_ADD100|32_  & ~new_n1104_;
  assign s33 = ~new_n1106_ & ~new_n1108_;
  assign \new_ADD100|33_  = new_n1100_ | new_n1106_;
  assign new_n1112_ = a34 & b34;
  assign new_n1114_ = ~a34 & ~b34;
  assign new_n1116_ = ~new_n1112_ & ~new_n1114_;
  assign new_n1118_ = \new_ADD100|33_  & new_n1116_;
  assign new_n1120_ = ~\new_ADD100|33_  & ~new_n1116_;
  assign s34 = ~new_n1118_ & ~new_n1120_;
  assign \new_ADD100|34_  = new_n1112_ | new_n1118_;
  assign new_n1124_ = a35 & b35;
  assign new_n1126_ = ~a35 & ~b35;
  assign new_n1128_ = ~new_n1124_ & ~new_n1126_;
  assign new_n1130_ = \new_ADD100|34_  & new_n1128_;
  assign new_n1132_ = ~\new_ADD100|34_  & ~new_n1128_;
  assign s35 = ~new_n1130_ & ~new_n1132_;
  assign \new_ADD100|35_  = new_n1124_ | new_n1130_;
  assign new_n1136_ = a36 & b36;
  assign new_n1138_ = ~a36 & ~b36;
  assign new_n1140_ = ~new_n1136_ & ~new_n1138_;
  assign new_n1142_ = \new_ADD100|35_  & new_n1140_;
  assign new_n1144_ = ~\new_ADD100|35_  & ~new_n1140_;
  assign s36 = ~new_n1142_ & ~new_n1144_;
  assign \new_ADD100|36_  = new_n1136_ | new_n1142_;
  assign new_n1148_ = a37 & b37;
  assign new_n1150_ = ~a37 & ~b37;
  assign new_n1152_ = ~new_n1148_ & ~new_n1150_;
  assign new_n1154_ = \new_ADD100|36_  & new_n1152_;
  assign new_n1156_ = ~\new_ADD100|36_  & ~new_n1152_;
  assign s37 = ~new_n1154_ & ~new_n1156_;
  assign \new_ADD100|37_  = new_n1148_ | new_n1154_;
  assign new_n1160_ = a38 & b38;
  assign new_n1162_ = ~a38 & ~b38;
  assign new_n1164_ = ~new_n1160_ & ~new_n1162_;
  assign new_n1166_ = \new_ADD100|37_  & new_n1164_;
  assign new_n1168_ = ~\new_ADD100|37_  & ~new_n1164_;
  assign s38 = ~new_n1166_ & ~new_n1168_;
  assign \new_ADD100|38_  = new_n1160_ | new_n1166_;
  assign new_n1172_ = a39 & b39;
  assign new_n1174_ = ~a39 & ~b39;
  assign new_n1176_ = ~new_n1172_ & ~new_n1174_;
  assign new_n1178_ = \new_ADD100|38_  & new_n1176_;
  assign new_n1180_ = ~\new_ADD100|38_  & ~new_n1176_;
  assign s39 = ~new_n1178_ & ~new_n1180_;
  assign \new_ADD100|39_  = new_n1172_ | new_n1178_;
  assign new_n1184_ = a40 & b40;
  assign new_n1186_ = ~a40 & ~b40;
  assign new_n1188_ = ~new_n1184_ & ~new_n1186_;
  assign new_n1190_ = \new_ADD100|39_  & new_n1188_;
  assign new_n1192_ = ~\new_ADD100|39_  & ~new_n1188_;
  assign s40 = ~new_n1190_ & ~new_n1192_;
  assign \new_ADD100|40_  = new_n1184_ | new_n1190_;
  assign new_n1196_ = a41 & b41;
  assign new_n1198_ = ~a41 & ~b41;
  assign new_n1200_ = ~new_n1196_ & ~new_n1198_;
  assign new_n1202_ = \new_ADD100|40_  & new_n1200_;
  assign new_n1204_ = ~\new_ADD100|40_  & ~new_n1200_;
  assign s41 = ~new_n1202_ & ~new_n1204_;
  assign \new_ADD100|41_  = new_n1196_ | new_n1202_;
  assign new_n1208_ = a42 & b42;
  assign new_n1210_ = ~a42 & ~b42;
  assign new_n1212_ = ~new_n1208_ & ~new_n1210_;
  assign new_n1214_ = \new_ADD100|41_  & new_n1212_;
  assign new_n1216_ = ~\new_ADD100|41_  & ~new_n1212_;
  assign s42 = ~new_n1214_ & ~new_n1216_;
  assign \new_ADD100|42_  = new_n1208_ | new_n1214_;
  assign new_n1220_ = a43 & b43;
  assign new_n1222_ = ~a43 & ~b43;
  assign new_n1224_ = ~new_n1220_ & ~new_n1222_;
  assign new_n1226_ = \new_ADD100|42_  & new_n1224_;
  assign new_n1228_ = ~\new_ADD100|42_  & ~new_n1224_;
  assign s43 = ~new_n1226_ & ~new_n1228_;
  assign \new_ADD100|43_  = new_n1220_ | new_n1226_;
  assign new_n1232_ = a44 & b44;
  assign new_n1234_ = ~a44 & ~b44;
  assign new_n1236_ = ~new_n1232_ & ~new_n1234_;
  assign new_n1238_ = \new_ADD100|43_  & new_n1236_;
  assign new_n1240_ = ~\new_ADD100|43_  & ~new_n1236_;
  assign s44 = ~new_n1238_ & ~new_n1240_;
  assign \new_ADD100|44_  = new_n1232_ | new_n1238_;
  assign new_n1244_ = a45 & b45;
  assign new_n1246_ = ~a45 & ~b45;
  assign new_n1248_ = ~new_n1244_ & ~new_n1246_;
  assign new_n1250_ = \new_ADD100|44_  & new_n1248_;
  assign new_n1252_ = ~\new_ADD100|44_  & ~new_n1248_;
  assign s45 = ~new_n1250_ & ~new_n1252_;
  assign \new_ADD100|45_  = new_n1244_ | new_n1250_;
  assign new_n1256_ = a46 & b46;
  assign new_n1258_ = ~a46 & ~b46;
  assign new_n1260_ = ~new_n1256_ & ~new_n1258_;
  assign new_n1262_ = \new_ADD100|45_  & new_n1260_;
  assign new_n1264_ = ~\new_ADD100|45_  & ~new_n1260_;
  assign s46 = ~new_n1262_ & ~new_n1264_;
  assign \new_ADD100|46_  = new_n1256_ | new_n1262_;
  assign new_n1268_ = a47 & b47;
  assign new_n1270_ = ~a47 & ~b47;
  assign new_n1272_ = ~new_n1268_ & ~new_n1270_;
  assign new_n1274_ = \new_ADD100|46_  & new_n1272_;
  assign new_n1276_ = ~\new_ADD100|46_  & ~new_n1272_;
  assign s47 = ~new_n1274_ & ~new_n1276_;
  assign \new_ADD100|47_  = new_n1268_ | new_n1274_;
  assign new_n1280_ = a48 & b48;
  assign new_n1282_ = ~a48 & ~b48;
  assign new_n1284_ = ~new_n1280_ & ~new_n1282_;
  assign new_n1286_ = \new_ADD100|47_  & new_n1284_;
  assign new_n1288_ = ~\new_ADD100|47_  & ~new_n1284_;
  assign s48 = ~new_n1286_ & ~new_n1288_;
  assign \new_ADD100|48_  = new_n1280_ | new_n1286_;
  assign new_n1292_ = a49 & b49;
  assign new_n1294_ = ~a49 & ~b49;
  assign new_n1296_ = ~new_n1292_ & ~new_n1294_;
  assign new_n1298_ = \new_ADD100|48_  & new_n1296_;
  assign new_n1300_ = ~\new_ADD100|48_  & ~new_n1296_;
  assign s49 = ~new_n1298_ & ~new_n1300_;
  assign \new_ADD100|49_  = new_n1292_ | new_n1298_;
  assign new_n1304_ = a50 & b50;
  assign new_n1306_ = ~a50 & ~b50;
  assign new_n1308_ = ~new_n1304_ & ~new_n1306_;
  assign new_n1310_ = \new_ADD100|49_  & new_n1308_;
  assign new_n1312_ = ~\new_ADD100|49_  & ~new_n1308_;
  assign s50 = ~new_n1310_ & ~new_n1312_;
  assign \new_ADD100|50_  = new_n1304_ | new_n1310_;
  assign new_n1316_ = a51 & b51;
  assign new_n1318_ = ~a51 & ~b51;
  assign new_n1320_ = ~new_n1316_ & ~new_n1318_;
  assign new_n1322_ = \new_ADD100|50_  & new_n1320_;
  assign new_n1324_ = ~\new_ADD100|50_  & ~new_n1320_;
  assign s51 = ~new_n1322_ & ~new_n1324_;
  assign \new_ADD100|51_  = new_n1316_ | new_n1322_;
  assign new_n1328_ = a52 & b52;
  assign new_n1330_ = ~a52 & ~b52;
  assign new_n1332_ = ~new_n1328_ & ~new_n1330_;
  assign new_n1334_ = \new_ADD100|51_  & new_n1332_;
  assign new_n1336_ = ~\new_ADD100|51_  & ~new_n1332_;
  assign s52 = ~new_n1334_ & ~new_n1336_;
  assign \new_ADD100|52_  = new_n1328_ | new_n1334_;
  assign new_n1340_ = a53 & b53;
  assign new_n1342_ = ~a53 & ~b53;
  assign new_n1344_ = ~new_n1340_ & ~new_n1342_;
  assign new_n1346_ = \new_ADD100|52_  & new_n1344_;
  assign new_n1348_ = ~\new_ADD100|52_  & ~new_n1344_;
  assign s53 = ~new_n1346_ & ~new_n1348_;
  assign \new_ADD100|53_  = new_n1340_ | new_n1346_;
  assign new_n1352_ = a54 & b54;
  assign new_n1354_ = ~a54 & ~b54;
  assign new_n1356_ = ~new_n1352_ & ~new_n1354_;
  assign new_n1358_ = \new_ADD100|53_  & new_n1356_;
  assign new_n1360_ = ~\new_ADD100|53_  & ~new_n1356_;
  assign s54 = ~new_n1358_ & ~new_n1360_;
  assign \new_ADD100|54_  = new_n1352_ | new_n1358_;
  assign new_n1364_ = a55 & b55;
  assign new_n1366_ = ~a55 & ~b55;
  assign new_n1368_ = ~new_n1364_ & ~new_n1366_;
  assign new_n1370_ = \new_ADD100|54_  & new_n1368_;
  assign new_n1372_ = ~\new_ADD100|54_  & ~new_n1368_;
  assign s55 = ~new_n1370_ & ~new_n1372_;
  assign \new_ADD100|55_  = new_n1364_ | new_n1370_;
  assign new_n1376_ = a56 & b56;
  assign new_n1378_ = ~a56 & ~b56;
  assign new_n1380_ = ~new_n1376_ & ~new_n1378_;
  assign new_n1382_ = \new_ADD100|55_  & new_n1380_;
  assign new_n1384_ = ~\new_ADD100|55_  & ~new_n1380_;
  assign s56 = ~new_n1382_ & ~new_n1384_;
  assign \new_ADD100|56_  = new_n1376_ | new_n1382_;
  assign new_n1388_ = a57 & b57;
  assign new_n1390_ = ~a57 & ~b57;
  assign new_n1392_ = ~new_n1388_ & ~new_n1390_;
  assign new_n1394_ = \new_ADD100|56_  & new_n1392_;
  assign new_n1396_ = ~\new_ADD100|56_  & ~new_n1392_;
  assign s57 = ~new_n1394_ & ~new_n1396_;
  assign \new_ADD100|57_  = new_n1388_ | new_n1394_;
  assign new_n1400_ = a58 & b58;
  assign new_n1402_ = ~a58 & ~b58;
  assign new_n1404_ = ~new_n1400_ & ~new_n1402_;
  assign new_n1406_ = \new_ADD100|57_  & new_n1404_;
  assign new_n1408_ = ~\new_ADD100|57_  & ~new_n1404_;
  assign s58 = ~new_n1406_ & ~new_n1408_;
  assign \new_ADD100|58_  = new_n1400_ | new_n1406_;
  assign new_n1412_ = a59 & b59;
  assign new_n1414_ = ~a59 & ~b59;
  assign new_n1416_ = ~new_n1412_ & ~new_n1414_;
  assign new_n1418_ = \new_ADD100|58_  & new_n1416_;
  assign new_n1420_ = ~\new_ADD100|58_  & ~new_n1416_;
  assign s59 = ~new_n1418_ & ~new_n1420_;
  assign \new_ADD100|59_  = new_n1412_ | new_n1418_;
  assign new_n1424_ = a60 & b60;
  assign new_n1426_ = ~a60 & ~b60;
  assign new_n1428_ = ~new_n1424_ & ~new_n1426_;
  assign new_n1430_ = \new_ADD100|59_  & new_n1428_;
  assign new_n1432_ = ~\new_ADD100|59_  & ~new_n1428_;
  assign s60 = ~new_n1430_ & ~new_n1432_;
  assign \new_ADD100|60_  = new_n1424_ | new_n1430_;
  assign new_n1436_ = a61 & b61;
  assign new_n1438_ = ~a61 & ~b61;
  assign new_n1440_ = ~new_n1436_ & ~new_n1438_;
  assign new_n1442_ = \new_ADD100|60_  & new_n1440_;
  assign new_n1444_ = ~\new_ADD100|60_  & ~new_n1440_;
  assign s61 = ~new_n1442_ & ~new_n1444_;
  assign \new_ADD100|61_  = new_n1436_ | new_n1442_;
  assign new_n1448_ = a62 & b62;
  assign new_n1450_ = ~a62 & ~b62;
  assign new_n1452_ = ~new_n1448_ & ~new_n1450_;
  assign new_n1454_ = \new_ADD100|61_  & new_n1452_;
  assign new_n1456_ = ~\new_ADD100|61_  & ~new_n1452_;
  assign s62 = ~new_n1454_ & ~new_n1456_;
  assign \new_ADD100|62_  = new_n1448_ | new_n1454_;
  assign new_n1460_ = a63 & b63;
  assign new_n1462_ = ~a63 & ~b63;
  assign new_n1464_ = ~new_n1460_ & ~new_n1462_;
  assign new_n1466_ = \new_ADD100|62_  & new_n1464_;
  assign new_n1468_ = ~\new_ADD100|62_  & ~new_n1464_;
  assign s63 = ~new_n1466_ & ~new_n1468_;
  assign \new_ADD100|63_  = new_n1460_ | new_n1466_;
  assign new_n1472_ = a64 & b64;
  assign new_n1474_ = ~a64 & ~b64;
  assign new_n1476_ = ~new_n1472_ & ~new_n1474_;
  assign new_n1478_ = \new_ADD100|63_  & new_n1476_;
  assign new_n1480_ = ~\new_ADD100|63_  & ~new_n1476_;
  assign s64 = ~new_n1478_ & ~new_n1480_;
  assign \new_ADD100|64_  = new_n1472_ | new_n1478_;
  assign new_n1484_ = a65 & b65;
  assign new_n1486_ = ~a65 & ~b65;
  assign new_n1488_ = ~new_n1484_ & ~new_n1486_;
  assign new_n1490_ = \new_ADD100|64_  & new_n1488_;
  assign new_n1492_ = ~\new_ADD100|64_  & ~new_n1488_;
  assign s65 = ~new_n1490_ & ~new_n1492_;
  assign \new_ADD100|65_  = new_n1484_ | new_n1490_;
  assign new_n1496_ = a66 & b66;
  assign new_n1498_ = ~a66 & ~b66;
  assign new_n1500_ = ~new_n1496_ & ~new_n1498_;
  assign new_n1502_ = \new_ADD100|65_  & new_n1500_;
  assign new_n1504_ = ~\new_ADD100|65_  & ~new_n1500_;
  assign s66 = ~new_n1502_ & ~new_n1504_;
  assign \new_ADD100|66_  = new_n1496_ | new_n1502_;
  assign new_n1508_ = a67 & b67;
  assign new_n1510_ = ~a67 & ~b67;
  assign new_n1512_ = ~new_n1508_ & ~new_n1510_;
  assign new_n1514_ = \new_ADD100|66_  & new_n1512_;
  assign new_n1516_ = ~\new_ADD100|66_  & ~new_n1512_;
  assign s67 = ~new_n1514_ & ~new_n1516_;
  assign \new_ADD100|67_  = new_n1508_ | new_n1514_;
  assign new_n1520_ = a68 & b68;
  assign new_n1522_ = ~a68 & ~b68;
  assign new_n1524_ = ~new_n1520_ & ~new_n1522_;
  assign new_n1526_ = \new_ADD100|67_  & new_n1524_;
  assign new_n1528_ = ~\new_ADD100|67_  & ~new_n1524_;
  assign s68 = ~new_n1526_ & ~new_n1528_;
  assign \new_ADD100|68_  = new_n1520_ | new_n1526_;
  assign new_n1532_ = a69 & b69;
  assign new_n1534_ = ~a69 & ~b69;
  assign new_n1536_ = ~new_n1532_ & ~new_n1534_;
  assign new_n1538_ = \new_ADD100|68_  & new_n1536_;
  assign new_n1540_ = ~\new_ADD100|68_  & ~new_n1536_;
  assign s69 = ~new_n1538_ & ~new_n1540_;
  assign \new_ADD100|69_  = new_n1532_ | new_n1538_;
  assign new_n1544_ = a70 & b70;
  assign new_n1546_ = ~a70 & ~b70;
  assign new_n1548_ = ~new_n1544_ & ~new_n1546_;
  assign new_n1550_ = \new_ADD100|69_  & new_n1548_;
  assign new_n1552_ = ~\new_ADD100|69_  & ~new_n1548_;
  assign s70 = ~new_n1550_ & ~new_n1552_;
  assign \new_ADD100|70_  = new_n1544_ | new_n1550_;
  assign new_n1556_ = a71 & b71;
  assign new_n1558_ = ~a71 & ~b71;
  assign new_n1560_ = ~new_n1556_ & ~new_n1558_;
  assign new_n1562_ = \new_ADD100|70_  & new_n1560_;
  assign new_n1564_ = ~\new_ADD100|70_  & ~new_n1560_;
  assign s71 = ~new_n1562_ & ~new_n1564_;
  assign \new_ADD100|71_  = new_n1556_ | new_n1562_;
  assign new_n1568_ = a72 & b72;
  assign new_n1570_ = ~a72 & ~b72;
  assign new_n1572_ = ~new_n1568_ & ~new_n1570_;
  assign new_n1574_ = \new_ADD100|71_  & new_n1572_;
  assign new_n1576_ = ~\new_ADD100|71_  & ~new_n1572_;
  assign s72 = ~new_n1574_ & ~new_n1576_;
  assign \new_ADD100|72_  = new_n1568_ | new_n1574_;
  assign new_n1580_ = a73 & b73;
  assign new_n1582_ = ~a73 & ~b73;
  assign new_n1584_ = ~new_n1580_ & ~new_n1582_;
  assign new_n1586_ = \new_ADD100|72_  & new_n1584_;
  assign new_n1588_ = ~\new_ADD100|72_  & ~new_n1584_;
  assign s73 = ~new_n1586_ & ~new_n1588_;
  assign \new_ADD100|73_  = new_n1580_ | new_n1586_;
  assign new_n1592_ = a74 & b74;
  assign new_n1594_ = ~a74 & ~b74;
  assign new_n1596_ = ~new_n1592_ & ~new_n1594_;
  assign new_n1598_ = \new_ADD100|73_  & new_n1596_;
  assign new_n1600_ = ~\new_ADD100|73_  & ~new_n1596_;
  assign s74 = ~new_n1598_ & ~new_n1600_;
  assign \new_ADD100|74_  = new_n1592_ | new_n1598_;
  assign new_n1604_ = a75 & b75;
  assign new_n1606_ = ~a75 & ~b75;
  assign new_n1608_ = ~new_n1604_ & ~new_n1606_;
  assign new_n1610_ = \new_ADD100|74_  & new_n1608_;
  assign new_n1612_ = ~\new_ADD100|74_  & ~new_n1608_;
  assign s75 = ~new_n1610_ & ~new_n1612_;
  assign \new_ADD100|75_  = new_n1604_ | new_n1610_;
  assign new_n1616_ = a76 & b76;
  assign new_n1618_ = ~a76 & ~b76;
  assign new_n1620_ = ~new_n1616_ & ~new_n1618_;
  assign new_n1622_ = \new_ADD100|75_  & new_n1620_;
  assign new_n1624_ = ~\new_ADD100|75_  & ~new_n1620_;
  assign s76 = ~new_n1622_ & ~new_n1624_;
  assign \new_ADD100|76_  = new_n1616_ | new_n1622_;
  assign new_n1628_ = a77 & b77;
  assign new_n1630_ = ~a77 & ~b77;
  assign new_n1632_ = ~new_n1628_ & ~new_n1630_;
  assign new_n1634_ = \new_ADD100|76_  & new_n1632_;
  assign new_n1636_ = ~\new_ADD100|76_  & ~new_n1632_;
  assign s77 = ~new_n1634_ & ~new_n1636_;
  assign \new_ADD100|77_  = new_n1628_ | new_n1634_;
  assign new_n1640_ = a78 & b78;
  assign new_n1642_ = ~a78 & ~b78;
  assign new_n1644_ = ~new_n1640_ & ~new_n1642_;
  assign new_n1646_ = \new_ADD100|77_  & new_n1644_;
  assign new_n1648_ = ~\new_ADD100|77_  & ~new_n1644_;
  assign s78 = ~new_n1646_ & ~new_n1648_;
  assign \new_ADD100|78_  = new_n1640_ | new_n1646_;
  assign new_n1652_ = a79 & b79;
  assign new_n1654_ = ~a79 & ~b79;
  assign new_n1656_ = ~new_n1652_ & ~new_n1654_;
  assign new_n1658_ = \new_ADD100|78_  & new_n1656_;
  assign new_n1660_ = ~\new_ADD100|78_  & ~new_n1656_;
  assign s79 = ~new_n1658_ & ~new_n1660_;
  assign \new_ADD100|79_  = new_n1652_ | new_n1658_;
  assign new_n1664_ = a80 & b80;
  assign new_n1666_ = ~a80 & ~b80;
  assign new_n1668_ = ~new_n1664_ & ~new_n1666_;
  assign new_n1670_ = \new_ADD100|79_  & new_n1668_;
  assign new_n1672_ = ~\new_ADD100|79_  & ~new_n1668_;
  assign s80 = ~new_n1670_ & ~new_n1672_;
  assign \new_ADD100|80_  = new_n1664_ | new_n1670_;
  assign new_n1676_ = a81 & b81;
  assign new_n1678_ = ~a81 & ~b81;
  assign new_n1680_ = ~new_n1676_ & ~new_n1678_;
  assign new_n1682_ = \new_ADD100|80_  & new_n1680_;
  assign new_n1684_ = ~\new_ADD100|80_  & ~new_n1680_;
  assign s81 = ~new_n1682_ & ~new_n1684_;
  assign \new_ADD100|81_  = new_n1676_ | new_n1682_;
  assign new_n1688_ = a82 & b82;
  assign new_n1690_ = ~a82 & ~b82;
  assign new_n1692_ = ~new_n1688_ & ~new_n1690_;
  assign new_n1694_ = \new_ADD100|81_  & new_n1692_;
  assign new_n1696_ = ~\new_ADD100|81_  & ~new_n1692_;
  assign s82 = ~new_n1694_ & ~new_n1696_;
  assign \new_ADD100|82_  = new_n1688_ | new_n1694_;
  assign new_n1700_ = a83 & b83;
  assign new_n1702_ = ~a83 & ~b83;
  assign new_n1704_ = ~new_n1700_ & ~new_n1702_;
  assign new_n1706_ = \new_ADD100|82_  & new_n1704_;
  assign new_n1708_ = ~\new_ADD100|82_  & ~new_n1704_;
  assign s83 = ~new_n1706_ & ~new_n1708_;
  assign \new_ADD100|83_  = new_n1700_ | new_n1706_;
  assign new_n1712_ = a84 & b84;
  assign new_n1714_ = ~a84 & ~b84;
  assign new_n1716_ = ~new_n1712_ & ~new_n1714_;
  assign new_n1718_ = \new_ADD100|83_  & new_n1716_;
  assign new_n1720_ = ~\new_ADD100|83_  & ~new_n1716_;
  assign s84 = ~new_n1718_ & ~new_n1720_;
  assign \new_ADD100|84_  = new_n1712_ | new_n1718_;
  assign new_n1724_ = a85 & b85;
  assign new_n1726_ = ~a85 & ~b85;
  assign new_n1728_ = ~new_n1724_ & ~new_n1726_;
  assign new_n1730_ = \new_ADD100|84_  & new_n1728_;
  assign new_n1732_ = ~\new_ADD100|84_  & ~new_n1728_;
  assign s85 = ~new_n1730_ & ~new_n1732_;
  assign \new_ADD100|85_  = new_n1724_ | new_n1730_;
  assign new_n1736_ = a86 & b86;
  assign new_n1738_ = ~a86 & ~b86;
  assign new_n1740_ = ~new_n1736_ & ~new_n1738_;
  assign new_n1742_ = \new_ADD100|85_  & new_n1740_;
  assign new_n1744_ = ~\new_ADD100|85_  & ~new_n1740_;
  assign s86 = ~new_n1742_ & ~new_n1744_;
  assign \new_ADD100|86_  = new_n1736_ | new_n1742_;
  assign new_n1748_ = a87 & b87;
  assign new_n1750_ = ~a87 & ~b87;
  assign new_n1752_ = ~new_n1748_ & ~new_n1750_;
  assign new_n1754_ = \new_ADD100|86_  & new_n1752_;
  assign new_n1756_ = ~\new_ADD100|86_  & ~new_n1752_;
  assign s87 = ~new_n1754_ & ~new_n1756_;
  assign \new_ADD100|87_  = new_n1748_ | new_n1754_;
  assign new_n1760_ = a88 & b88;
  assign new_n1762_ = ~a88 & ~b88;
  assign new_n1764_ = ~new_n1760_ & ~new_n1762_;
  assign new_n1766_ = \new_ADD100|87_  & new_n1764_;
  assign new_n1768_ = ~\new_ADD100|87_  & ~new_n1764_;
  assign s88 = ~new_n1766_ & ~new_n1768_;
  assign \new_ADD100|88_  = new_n1760_ | new_n1766_;
  assign new_n1772_ = a89 & b89;
  assign new_n1774_ = ~a89 & ~b89;
  assign new_n1776_ = ~new_n1772_ & ~new_n1774_;
  assign new_n1778_ = \new_ADD100|88_  & new_n1776_;
  assign new_n1780_ = ~\new_ADD100|88_  & ~new_n1776_;
  assign s89 = ~new_n1778_ & ~new_n1780_;
  assign \new_ADD100|89_  = new_n1772_ | new_n1778_;
  assign new_n1784_ = a90 & b90;
  assign new_n1786_ = ~a90 & ~b90;
  assign new_n1788_ = ~new_n1784_ & ~new_n1786_;
  assign new_n1790_ = \new_ADD100|89_  & new_n1788_;
  assign new_n1792_ = ~\new_ADD100|89_  & ~new_n1788_;
  assign s90 = ~new_n1790_ & ~new_n1792_;
  assign \new_ADD100|90_  = new_n1784_ | new_n1790_;
  assign new_n1796_ = a91 & b91;
  assign new_n1798_ = ~a91 & ~b91;
  assign new_n1800_ = ~new_n1796_ & ~new_n1798_;
  assign new_n1802_ = \new_ADD100|90_  & new_n1800_;
  assign new_n1804_ = ~\new_ADD100|90_  & ~new_n1800_;
  assign s91 = ~new_n1802_ & ~new_n1804_;
  assign \new_ADD100|91_  = new_n1796_ | new_n1802_;
  assign new_n1808_ = a92 & b92;
  assign new_n1810_ = ~a92 & ~b92;
  assign new_n1812_ = ~new_n1808_ & ~new_n1810_;
  assign new_n1814_ = \new_ADD100|91_  & new_n1812_;
  assign new_n1816_ = ~\new_ADD100|91_  & ~new_n1812_;
  assign s92 = ~new_n1814_ & ~new_n1816_;
  assign \new_ADD100|92_  = new_n1808_ | new_n1814_;
  assign new_n1820_ = a93 & b93;
  assign new_n1822_ = ~a93 & ~b93;
  assign new_n1824_ = ~new_n1820_ & ~new_n1822_;
  assign new_n1826_ = \new_ADD100|92_  & new_n1824_;
  assign new_n1828_ = ~\new_ADD100|92_  & ~new_n1824_;
  assign s93 = ~new_n1826_ & ~new_n1828_;
  assign \new_ADD100|93_  = new_n1820_ | new_n1826_;
  assign new_n1832_ = a94 & b94;
  assign new_n1834_ = ~a94 & ~b94;
  assign new_n1836_ = ~new_n1832_ & ~new_n1834_;
  assign new_n1838_ = \new_ADD100|93_  & new_n1836_;
  assign new_n1840_ = ~\new_ADD100|93_  & ~new_n1836_;
  assign s94 = ~new_n1838_ & ~new_n1840_;
  assign \new_ADD100|94_  = new_n1832_ | new_n1838_;
  assign new_n1844_ = a95 & b95;
  assign new_n1846_ = ~a95 & ~b95;
  assign new_n1848_ = ~new_n1844_ & ~new_n1846_;
  assign new_n1850_ = \new_ADD100|94_  & new_n1848_;
  assign new_n1852_ = ~\new_ADD100|94_  & ~new_n1848_;
  assign s95 = ~new_n1850_ & ~new_n1852_;
  assign \new_ADD100|95_  = new_n1844_ | new_n1850_;
  assign new_n1856_ = a96 & b96;
  assign new_n1858_ = ~a96 & ~b96;
  assign new_n1860_ = ~new_n1856_ & ~new_n1858_;
  assign new_n1862_ = \new_ADD100|95_  & new_n1860_;
  assign new_n1864_ = ~\new_ADD100|95_  & ~new_n1860_;
  assign s96 = ~new_n1862_ & ~new_n1864_;
  assign \new_ADD100|96_  = new_n1856_ | new_n1862_;
  assign new_n1868_ = a97 & b97;
  assign new_n1870_ = ~a97 & ~b97;
  assign new_n1872_ = ~new_n1868_ & ~new_n1870_;
  assign new_n1874_ = \new_ADD100|96_  & new_n1872_;
  assign new_n1876_ = ~\new_ADD100|96_  & ~new_n1872_;
  assign s97 = ~new_n1874_ & ~new_n1876_;
  assign \new_ADD100|97_  = new_n1868_ | new_n1874_;
  assign new_n1880_ = a98 & b98;
  assign new_n1882_ = ~a98 & ~b98;
  assign new_n1884_ = ~new_n1880_ & ~new_n1882_;
  assign new_n1886_ = \new_ADD100|97_  & new_n1884_;
  assign new_n1888_ = ~\new_ADD100|97_  & ~new_n1884_;
  assign s98 = ~new_n1886_ & ~new_n1888_;
  assign \new_ADD100|98_  = new_n1880_ | new_n1886_;
  assign new_n1892_ = a99 & b99;
  assign new_n1894_ = ~a99 & ~b99;
  assign new_n1896_ = ~new_n1892_ & ~new_n1894_;
  assign new_n1898_ = \new_ADD100|98_  & new_n1896_;
  assign new_n1900_ = ~\new_ADD100|98_  & ~new_n1896_;
  assign s99 = ~new_n1898_ & ~new_n1900_;
  assign s100 = new_n1892_ | new_n1898_;
endmodule


